module test_16( pi0, pi1, pi2, pi3, pi4, po0 );
  input pi0, pi1, pi2, pi3, pi4;
  output po0;
  wire w1;
  wire tmp0;
  assign tmp0 = 1'b1;
  wire tmp1;
  assign tmp1 = pi0;
  wire tmp2;
  assign tmp2 = pi1;
  wire tmp3;
  assign tmp3 = (tmp0 & tmp1) | (tmp0 & tmp2) | (tmp1 & tmp2);
  wire tmp4;
  assign tmp4 = pi0;
  wire tmp5;
  assign tmp5 = 1'b1;
  wire tmp6;
  assign tmp6 = 1'b1;
  wire tmp7;
  assign tmp7 = (tmp4 & tmp5) | (tmp4 & tmp6) | (tmp5 & tmp6);
  wire tmp8;
  assign tmp8 = pi1;
  wire tmp9;
  assign tmp9 = 1'b1;
  wire tmp10;
  assign tmp10 = 1'b0;
  wire tmp11;
  assign tmp11 = (tmp8 & tmp9) | (tmp8 & tmp10) | (tmp9 & tmp10);
  wire tmp12;
  assign tmp12 = (tmp3 & tmp7) | (tmp3 & tmp11) | (tmp7 & tmp11);
  assign w1 = tmp12;
  wire tmp13;
  assign tmp13 = w1;
  wire tmp14;
  assign tmp14 = ~pi4;
  wire tmp15;
  assign tmp15 = 1'b0;
  wire tmp16;
  assign tmp16 = (tmp13 & tmp14) | (tmp13 & tmp15) | (tmp14 & tmp15);
  wire tmp17;
  assign tmp17 = ~pi4;
  wire tmp18;
  assign tmp18 = ~pi2;
  wire tmp19;
  assign tmp19 = 1'b0;
  wire tmp20;
  assign tmp20 = (tmp17 & tmp18) | (tmp17 & tmp19) | (tmp18 & tmp19);
  wire tmp21;
  assign tmp21 = 1'b0;
  wire tmp22;
  assign tmp22 = 1'b0;
  wire tmp23;
  assign tmp23 = 1'b0;
  wire tmp24;
  assign tmp24 = (tmp21 & tmp22) | (tmp21 & tmp23) | (tmp22 & tmp23);
  wire tmp25;
  assign tmp25 = (tmp16 & tmp20) | (tmp16 & tmp24) | (tmp20 & tmp24);
  wire tmp26;
  assign tmp26 = ~pi4;
  wire tmp27;
  assign tmp27 = ~pi2;
  wire tmp28;
  assign tmp28 = 1'b0;
  wire tmp29;
  assign tmp29 = (tmp26 & tmp27) | (tmp26 & tmp28) | (tmp27 & tmp28);
  wire tmp30;
  assign tmp30 = ~pi2;
  wire tmp31;
  assign tmp31 = ~pi3;
  wire tmp32;
  assign tmp32 = 1'b0;
  wire tmp33;
  assign tmp33 = (tmp30 & tmp31) | (tmp30 & tmp32) | (tmp31 & tmp32);
  wire tmp34;
  assign tmp34 = 1'b0;
  wire tmp35;
  assign tmp35 = 1'b0;
  wire tmp36;
  assign tmp36 = 1'b0;
  wire tmp37;
  assign tmp37 = (tmp34 & tmp35) | (tmp34 & tmp36) | (tmp35 & tmp36);
  wire tmp38;
  assign tmp38 = (tmp29 & tmp33) | (tmp29 & tmp37) | (tmp33 & tmp37);
  wire tmp39;
  assign tmp39 = 1'b0;
  wire tmp40;
  assign tmp40 = 1'b0;
  wire tmp41;
  assign tmp41 = 1'b0;
  wire tmp42;
  assign tmp42 = (tmp39 & tmp40) | (tmp39 & tmp41) | (tmp40 & tmp41);
  wire tmp43;
  assign tmp43 = 1'b0;
  wire tmp44;
  assign tmp44 = 1'b0;
  wire tmp45;
  assign tmp45 = 1'b0;
  wire tmp46;
  assign tmp46 = (tmp43 & tmp44) | (tmp43 & tmp45) | (tmp44 & tmp45);
  wire tmp47;
  assign tmp47 = 1'b0;
  wire tmp48;
  assign tmp48 = 1'b0;
  wire tmp49;
  assign tmp49 = 1'b0;
  wire tmp50;
  assign tmp50 = (tmp47 & tmp48) | (tmp47 & tmp49) | (tmp48 & tmp49);
  wire tmp51;
  assign tmp51 = (tmp42 & tmp46) | (tmp42 & tmp50) | (tmp46 & tmp50);
  wire tmp52;
  assign tmp52 = (tmp25 & tmp38) | (tmp25 & tmp51) | (tmp38 & tmp51);
  assign po0 = tmp52;
endmodule // test_16
