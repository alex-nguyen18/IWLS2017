module test_each( pi0, pi1, pi2, pi3, pi4, pi5, po0, po1, po2, po3, po4, po5 );
  input pi0, pi1, pi2, pi3, pi4, pi5;
  output po0, po1, po2, po3, po4, po5;
  wire w1;
  wire tmp0;
  assign tmp0 = pi2;
  wire tmp1;
  assign tmp1 = pi3;
  wire tmp2;
  assign tmp2 = 1'b0;
  wire tmp3;
  assign tmp3 = (tmp0 & tmp1) | (tmp0 & tmp2) | (tmp1 & tmp2);
  assign w1 = tmp3;
  wire tmp4;
  assign tmp4 = pi0;
  wire tmp5;
  assign tmp5 = pi1;
  wire tmp6;
  assign tmp6 = 1'b0;
  wire tmp7;
  assign tmp7 = (tmp4 & tmp5) | (tmp4 & tmp6) | (tmp5 & tmp6);
  assign po0 = tmp7;
  wire tmp8;
  assign tmp8 = 1'b1;
  wire tmp9;
  assign tmp9 = pi0;
  wire tmp10;
  assign tmp10 = pi1;
  wire tmp11;
  assign tmp11 = (tmp8 & tmp9) | (tmp8 & tmp10) | (tmp9 & tmp10);
  wire tmp12;
  assign tmp12 = pi0;
  wire tmp13;
  assign tmp13 = 1'b1;
  wire tmp14;
  assign tmp14 = 1'b1;
  wire tmp15;
  assign tmp15 = (tmp12 & tmp13) | (tmp12 & tmp14) | (tmp13 & tmp14);
  wire tmp16;
  assign tmp16 = pi1;
  wire tmp17;
  assign tmp17 = 1'b1;
  wire tmp18;
  assign tmp18 = 1'b0;
  wire tmp19;
  assign tmp19 = (tmp16 & tmp17) | (tmp16 & tmp18) | (tmp17 & tmp18);
  wire tmp20;
  assign tmp20 = (tmp11 & tmp15) | (tmp11 & tmp19) | (tmp15 & tmp19);
  assign po1 = tmp20;
  wire tmp21;
  assign tmp21 = pi0;
  wire tmp22;
  assign tmp22 = pi1;
  wire tmp23;
  assign tmp23 = 1'b0;
  wire tmp24;
  assign tmp24 = (tmp21 & tmp22) | (tmp21 & tmp23) | (tmp22 & tmp23);
  wire tmp25;
  assign tmp25 = pi1;
  wire tmp26;
  assign tmp26 = pi2;
  wire tmp27;
  assign tmp27 = 1'b0;
  wire tmp28;
  assign tmp28 = (tmp25 & tmp26) | (tmp25 & tmp27) | (tmp26 & tmp27);
  wire tmp29;
  assign tmp29 = 1'b0;
  wire tmp30;
  assign tmp30 = 1'b0;
  wire tmp31;
  assign tmp31 = 1'b0;
  wire tmp32;
  assign tmp32 = (tmp29 & tmp30) | (tmp29 & tmp31) | (tmp30 & tmp31);
  wire tmp33;
  assign tmp33 = (tmp24 & tmp28) | (tmp24 & tmp32) | (tmp28 & tmp32);
  wire tmp34;
  assign tmp34 = pi1;
  wire tmp35;
  assign tmp35 = pi2;
  wire tmp36;
  assign tmp36 = 1'b0;
  wire tmp37;
  assign tmp37 = (tmp34 & tmp35) | (tmp34 & tmp36) | (tmp35 & tmp36);
  wire tmp38;
  assign tmp38 = pi2;
  wire tmp39;
  assign tmp39 = pi3;
  wire tmp40;
  assign tmp40 = 1'b0;
  wire tmp41;
  assign tmp41 = (tmp38 & tmp39) | (tmp38 & tmp40) | (tmp39 & tmp40);
  wire tmp42;
  assign tmp42 = 1'b0;
  wire tmp43;
  assign tmp43 = 1'b0;
  wire tmp44;
  assign tmp44 = 1'b0;
  wire tmp45;
  assign tmp45 = (tmp42 & tmp43) | (tmp42 & tmp44) | (tmp43 & tmp44);
  wire tmp46;
  assign tmp46 = (tmp37 & tmp41) | (tmp37 & tmp45) | (tmp41 & tmp45);
  wire tmp47;
  assign tmp47 = 1'b0;
  wire tmp48;
  assign tmp48 = 1'b0;
  wire tmp49;
  assign tmp49 = 1'b0;
  wire tmp50;
  assign tmp50 = (tmp47 & tmp48) | (tmp47 & tmp49) | (tmp48 & tmp49);
  wire tmp51;
  assign tmp51 = 1'b0;
  wire tmp52;
  assign tmp52 = 1'b0;
  wire tmp53;
  assign tmp53 = 1'b0;
  wire tmp54;
  assign tmp54 = (tmp51 & tmp52) | (tmp51 & tmp53) | (tmp52 & tmp53);
  wire tmp55;
  assign tmp55 = 1'b0;
  wire tmp56;
  assign tmp56 = 1'b0;
  wire tmp57;
  assign tmp57 = 1'b0;
  wire tmp58;
  assign tmp58 = (tmp55 & tmp56) | (tmp55 & tmp57) | (tmp56 & tmp57);
  wire tmp59;
  assign tmp59 = (tmp50 & tmp54) | (tmp50 & tmp58) | (tmp54 & tmp58);
  wire tmp60;
  assign tmp60 = (tmp33 & tmp46) | (tmp33 & tmp59) | (tmp46 & tmp59);
  assign po2 = tmp60;
  wire tmp61;
  assign tmp61 = 1'b1;
  wire tmp62;
  assign tmp62 = 1'b1;
  wire tmp63;
  assign tmp63 = 1'b1;
  wire tmp64;
  assign tmp64 = (tmp61 & tmp62) | (tmp61 & tmp63) | (tmp62 & tmp63);
  wire tmp65;
  assign tmp65 = 1'b1;
  wire tmp66;
  assign tmp66 = 1'b1;
  wire tmp67;
  assign tmp67 = 1'b1;
  wire tmp68;
  assign tmp68 = (tmp65 & tmp66) | (tmp65 & tmp67) | (tmp66 & tmp67);
  wire tmp69;
  assign tmp69 = 1'b1;
  wire tmp70;
  assign tmp70 = 1'b1;
  wire tmp71;
  assign tmp71 = 1'b1;
  wire tmp72;
  assign tmp72 = (tmp69 & tmp70) | (tmp69 & tmp71) | (tmp70 & tmp71);
  wire tmp73;
  assign tmp73 = (tmp64 & tmp68) | (tmp64 & tmp72) | (tmp68 & tmp72);
  wire tmp74;
  assign tmp74 = 1'b1;
  wire tmp75;
  assign tmp75 = 1'b1;
  wire tmp76;
  assign tmp76 = 1'b1;
  wire tmp77;
  assign tmp77 = (tmp74 & tmp75) | (tmp74 & tmp76) | (tmp75 & tmp76);
  wire tmp78;
  assign tmp78 = 1'b1;
  wire tmp79;
  assign tmp79 = pi0;
  wire tmp80;
  assign tmp80 = pi1;
  wire tmp81;
  assign tmp81 = (tmp78 & tmp79) | (tmp78 & tmp80) | (tmp79 & tmp80);
  wire tmp82;
  assign tmp82 = 1'b1;
  wire tmp83;
  assign tmp83 = pi1;
  wire tmp84;
  assign tmp84 = pi4;
  wire tmp85;
  assign tmp85 = (tmp82 & tmp83) | (tmp82 & tmp84) | (tmp83 & tmp84);
  wire tmp86;
  assign tmp86 = (tmp77 & tmp81) | (tmp77 & tmp85) | (tmp81 & tmp85);
  wire tmp87;
  assign tmp87 = 1'b1;
  wire tmp88;
  assign tmp88 = 1'b1;
  wire tmp89;
  assign tmp89 = 1'b1;
  wire tmp90;
  assign tmp90 = (tmp87 & tmp88) | (tmp87 & tmp89) | (tmp88 & tmp89);
  wire tmp91;
  assign tmp91 = 1'b1;
  wire tmp92;
  assign tmp92 = pi1;
  wire tmp93;
  assign tmp93 = pi4;
  wire tmp94;
  assign tmp94 = (tmp91 & tmp92) | (tmp91 & tmp93) | (tmp92 & tmp93);
  wire tmp95;
  assign tmp95 = 1'b1;
  wire tmp96;
  assign tmp96 = pi4;
  wire tmp97;
  assign tmp97 = pi5;
  wire tmp98;
  assign tmp98 = (tmp95 & tmp96) | (tmp95 & tmp97) | (tmp96 & tmp97);
  wire tmp99;
  assign tmp99 = (tmp90 & tmp94) | (tmp90 & tmp98) | (tmp94 & tmp98);
  wire tmp100;
  assign tmp100 = (tmp73 & tmp86) | (tmp73 & tmp99) | (tmp86 & tmp99);
  wire tmp101;
  assign tmp101 = 1'b1;
  wire tmp102;
  assign tmp102 = 1'b1;
  wire tmp103;
  assign tmp103 = 1'b1;
  wire tmp104;
  assign tmp104 = (tmp101 & tmp102) | (tmp101 & tmp103) | (tmp102 & tmp103);
  wire tmp105;
  assign tmp105 = 1'b1;
  wire tmp106;
  assign tmp106 = pi0;
  wire tmp107;
  assign tmp107 = pi1;
  wire tmp108;
  assign tmp108 = (tmp105 & tmp106) | (tmp105 & tmp107) | (tmp106 & tmp107);
  wire tmp109;
  assign tmp109 = 1'b1;
  wire tmp110;
  assign tmp110 = pi1;
  wire tmp111;
  assign tmp111 = pi4;
  wire tmp112;
  assign tmp112 = (tmp109 & tmp110) | (tmp109 & tmp111) | (tmp110 & tmp111);
  wire tmp113;
  assign tmp113 = (tmp104 & tmp108) | (tmp104 & tmp112) | (tmp108 & tmp112);
  wire tmp114;
  assign tmp114 = 1'b1;
  wire tmp115;
  assign tmp115 = pi0;
  wire tmp116;
  assign tmp116 = pi1;
  wire tmp117;
  assign tmp117 = (tmp114 & tmp115) | (tmp114 & tmp116) | (tmp115 & tmp116);
  wire tmp118;
  assign tmp118 = pi0;
  wire tmp119;
  assign tmp119 = 1'b1;
  wire tmp120;
  assign tmp120 = 1'b1;
  wire tmp121;
  assign tmp121 = (tmp118 & tmp119) | (tmp118 & tmp120) | (tmp119 & tmp120);
  wire tmp122;
  assign tmp122 = pi1;
  wire tmp123;
  assign tmp123 = 1'b1;
  wire tmp124;
  assign tmp124 = 1'b1;
  wire tmp125;
  assign tmp125 = (tmp122 & tmp123) | (tmp122 & tmp124) | (tmp123 & tmp124);
  wire tmp126;
  assign tmp126 = (tmp117 & tmp121) | (tmp117 & tmp125) | (tmp121 & tmp125);
  wire tmp127;
  assign tmp127 = 1'b1;
  wire tmp128;
  assign tmp128 = pi1;
  wire tmp129;
  assign tmp129 = pi4;
  wire tmp130;
  assign tmp130 = (tmp127 & tmp128) | (tmp127 & tmp129) | (tmp128 & tmp129);
  wire tmp131;
  assign tmp131 = pi1;
  wire tmp132;
  assign tmp132 = 1'b1;
  wire tmp133;
  assign tmp133 = 1'b1;
  wire tmp134;
  assign tmp134 = (tmp131 & tmp132) | (tmp131 & tmp133) | (tmp132 & tmp133);
  wire tmp135;
  assign tmp135 = pi4;
  wire tmp136;
  assign tmp136 = 1'b1;
  wire tmp137;
  assign tmp137 = 1'b1;
  wire tmp138;
  assign tmp138 = (tmp135 & tmp136) | (tmp135 & tmp137) | (tmp136 & tmp137);
  wire tmp139;
  assign tmp139 = (tmp130 & tmp134) | (tmp130 & tmp138) | (tmp134 & tmp138);
  wire tmp140;
  assign tmp140 = (tmp113 & tmp126) | (tmp113 & tmp139) | (tmp126 & tmp139);
  wire tmp141;
  assign tmp141 = 1'b1;
  wire tmp142;
  assign tmp142 = 1'b1;
  wire tmp143;
  assign tmp143 = 1'b1;
  wire tmp144;
  assign tmp144 = (tmp141 & tmp142) | (tmp141 & tmp143) | (tmp142 & tmp143);
  wire tmp145;
  assign tmp145 = 1'b1;
  wire tmp146;
  assign tmp146 = pi1;
  wire tmp147;
  assign tmp147 = pi4;
  wire tmp148;
  assign tmp148 = (tmp145 & tmp146) | (tmp145 & tmp147) | (tmp146 & tmp147);
  wire tmp149;
  assign tmp149 = 1'b1;
  wire tmp150;
  assign tmp150 = pi4;
  wire tmp151;
  assign tmp151 = pi5;
  wire tmp152;
  assign tmp152 = (tmp149 & tmp150) | (tmp149 & tmp151) | (tmp150 & tmp151);
  wire tmp153;
  assign tmp153 = (tmp144 & tmp148) | (tmp144 & tmp152) | (tmp148 & tmp152);
  wire tmp154;
  assign tmp154 = 1'b1;
  wire tmp155;
  assign tmp155 = pi1;
  wire tmp156;
  assign tmp156 = pi4;
  wire tmp157;
  assign tmp157 = (tmp154 & tmp155) | (tmp154 & tmp156) | (tmp155 & tmp156);
  wire tmp158;
  assign tmp158 = pi1;
  wire tmp159;
  assign tmp159 = 1'b1;
  wire tmp160;
  assign tmp160 = 1'b1;
  wire tmp161;
  assign tmp161 = (tmp158 & tmp159) | (tmp158 & tmp160) | (tmp159 & tmp160);
  wire tmp162;
  assign tmp162 = pi4;
  wire tmp163;
  assign tmp163 = 1'b1;
  wire tmp164;
  assign tmp164 = 1'b1;
  wire tmp165;
  assign tmp165 = (tmp162 & tmp163) | (tmp162 & tmp164) | (tmp163 & tmp164);
  wire tmp166;
  assign tmp166 = (tmp157 & tmp161) | (tmp157 & tmp165) | (tmp161 & tmp165);
  wire tmp167;
  assign tmp167 = 1'b1;
  wire tmp168;
  assign tmp168 = pi4;
  wire tmp169;
  assign tmp169 = pi5;
  wire tmp170;
  assign tmp170 = (tmp167 & tmp168) | (tmp167 & tmp169) | (tmp168 & tmp169);
  wire tmp171;
  assign tmp171 = pi4;
  wire tmp172;
  assign tmp172 = 1'b1;
  wire tmp173;
  assign tmp173 = 1'b1;
  wire tmp174;
  assign tmp174 = (tmp171 & tmp172) | (tmp171 & tmp173) | (tmp172 & tmp173);
  wire tmp175;
  assign tmp175 = pi5;
  wire tmp176;
  assign tmp176 = 1'b1;
  wire tmp177;
  assign tmp177 = 1'b0;
  wire tmp178;
  assign tmp178 = (tmp175 & tmp176) | (tmp175 & tmp177) | (tmp176 & tmp177);
  wire tmp179;
  assign tmp179 = (tmp170 & tmp174) | (tmp170 & tmp178) | (tmp174 & tmp178);
  wire tmp180;
  assign tmp180 = (tmp153 & tmp166) | (tmp153 & tmp179) | (tmp166 & tmp179);
  wire tmp181;
  assign tmp181 = (tmp100 & tmp140) | (tmp100 & tmp180) | (tmp140 & tmp180);
  assign po3 = tmp181;
  wire tmp182;
  assign tmp182 = pi2;
  wire tmp183;
  assign tmp183 = pi3;
  wire tmp184;
  assign tmp184 = 1'b0;
  wire tmp185;
  assign tmp185 = (tmp182 & tmp183) | (tmp182 & tmp184) | (tmp183 & tmp184);
  wire tmp186;
  assign tmp186 = pi3;
  wire tmp187;
  assign tmp187 = 1'b1;
  wire tmp188;
  assign tmp188 = 1'b0;
  wire tmp189;
  assign tmp189 = (tmp186 & tmp187) | (tmp186 & tmp188) | (tmp187 & tmp188);
  wire tmp190;
  assign tmp190 = 1'b0;
  wire tmp191;
  assign tmp191 = 1'b0;
  wire tmp192;
  assign tmp192 = 1'b0;
  wire tmp193;
  assign tmp193 = (tmp190 & tmp191) | (tmp190 & tmp192) | (tmp191 & tmp192);
  wire tmp194;
  assign tmp194 = (tmp185 & tmp189) | (tmp185 & tmp193) | (tmp189 & tmp193);
  wire tmp195;
  assign tmp195 = pi3;
  wire tmp196;
  assign tmp196 = 1'b1;
  wire tmp197;
  assign tmp197 = 1'b0;
  wire tmp198;
  assign tmp198 = (tmp195 & tmp196) | (tmp195 & tmp197) | (tmp196 & tmp197);
  wire tmp199;
  assign tmp199 = 1'b1;
  wire tmp200;
  assign tmp200 = pi4;
  wire tmp201;
  assign tmp201 = pi5;
  wire tmp202;
  assign tmp202 = (tmp199 & tmp200) | (tmp199 & tmp201) | (tmp200 & tmp201);
  wire tmp203;
  assign tmp203 = 1'b0;
  wire tmp204;
  assign tmp204 = pi5;
  wire tmp205;
  assign tmp205 = 1'b0;
  wire tmp206;
  assign tmp206 = (tmp203 & tmp204) | (tmp203 & tmp205) | (tmp204 & tmp205);
  wire tmp207;
  assign tmp207 = (tmp198 & tmp202) | (tmp198 & tmp206) | (tmp202 & tmp206);
  wire tmp208;
  assign tmp208 = 1'b0;
  wire tmp209;
  assign tmp209 = 1'b0;
  wire tmp210;
  assign tmp210 = 1'b0;
  wire tmp211;
  assign tmp211 = (tmp208 & tmp209) | (tmp208 & tmp210) | (tmp209 & tmp210);
  wire tmp212;
  assign tmp212 = 1'b0;
  wire tmp213;
  assign tmp213 = pi5;
  wire tmp214;
  assign tmp214 = 1'b0;
  wire tmp215;
  assign tmp215 = (tmp212 & tmp213) | (tmp212 & tmp214) | (tmp213 & tmp214);
  wire tmp216;
  assign tmp216 = 1'b0;
  wire tmp217;
  assign tmp217 = 1'b0;
  wire tmp218;
  assign tmp218 = 1'b0;
  wire tmp219;
  assign tmp219 = (tmp216 & tmp217) | (tmp216 & tmp218) | (tmp217 & tmp218);
  wire tmp220;
  assign tmp220 = (tmp211 & tmp215) | (tmp211 & tmp219) | (tmp215 & tmp219);
  wire tmp221;
  assign tmp221 = (tmp194 & tmp207) | (tmp194 & tmp220) | (tmp207 & tmp220);
  wire tmp222;
  assign tmp222 = pi3;
  wire tmp223;
  assign tmp223 = 1'b1;
  wire tmp224;
  assign tmp224 = 1'b0;
  wire tmp225;
  assign tmp225 = (tmp222 & tmp223) | (tmp222 & tmp224) | (tmp223 & tmp224);
  wire tmp226;
  assign tmp226 = 1'b1;
  wire tmp227;
  assign tmp227 = pi4;
  wire tmp228;
  assign tmp228 = pi5;
  wire tmp229;
  assign tmp229 = (tmp226 & tmp227) | (tmp226 & tmp228) | (tmp227 & tmp228);
  wire tmp230;
  assign tmp230 = 1'b0;
  wire tmp231;
  assign tmp231 = pi5;
  wire tmp232;
  assign tmp232 = 1'b0;
  wire tmp233;
  assign tmp233 = (tmp230 & tmp231) | (tmp230 & tmp232) | (tmp231 & tmp232);
  wire tmp234;
  assign tmp234 = (tmp225 & tmp229) | (tmp225 & tmp233) | (tmp229 & tmp233);
  wire tmp235;
  assign tmp235 = 1'b1;
  wire tmp236;
  assign tmp236 = pi4;
  wire tmp237;
  assign tmp237 = pi5;
  wire tmp238;
  assign tmp238 = (tmp235 & tmp236) | (tmp235 & tmp237) | (tmp236 & tmp237);
  wire tmp239;
  assign tmp239 = pi4;
  wire tmp240;
  assign tmp240 = 1'b1;
  wire tmp241;
  assign tmp241 = 1'b1;
  wire tmp242;
  assign tmp242 = (tmp239 & tmp240) | (tmp239 & tmp241) | (tmp240 & tmp241);
  wire tmp243;
  assign tmp243 = pi5;
  wire tmp244;
  assign tmp244 = 1'b1;
  wire tmp245;
  assign tmp245 = 1'b0;
  wire tmp246;
  assign tmp246 = (tmp243 & tmp244) | (tmp243 & tmp245) | (tmp244 & tmp245);
  wire tmp247;
  assign tmp247 = (tmp238 & tmp242) | (tmp238 & tmp246) | (tmp242 & tmp246);
  wire tmp248;
  assign tmp248 = 1'b0;
  wire tmp249;
  assign tmp249 = pi5;
  wire tmp250;
  assign tmp250 = 1'b0;
  wire tmp251;
  assign tmp251 = (tmp248 & tmp249) | (tmp248 & tmp250) | (tmp249 & tmp250);
  wire tmp252;
  assign tmp252 = pi5;
  wire tmp253;
  assign tmp253 = 1'b1;
  wire tmp254;
  assign tmp254 = 1'b0;
  wire tmp255;
  assign tmp255 = (tmp252 & tmp253) | (tmp252 & tmp254) | (tmp253 & tmp254);
  wire tmp256;
  assign tmp256 = 1'b0;
  wire tmp257;
  assign tmp257 = 1'b0;
  wire tmp258;
  assign tmp258 = 1'b0;
  wire tmp259;
  assign tmp259 = (tmp256 & tmp257) | (tmp256 & tmp258) | (tmp257 & tmp258);
  wire tmp260;
  assign tmp260 = (tmp251 & tmp255) | (tmp251 & tmp259) | (tmp255 & tmp259);
  wire tmp261;
  assign tmp261 = (tmp234 & tmp247) | (tmp234 & tmp260) | (tmp247 & tmp260);
  wire tmp262;
  assign tmp262 = 1'b0;
  wire tmp263;
  assign tmp263 = 1'b0;
  wire tmp264;
  assign tmp264 = 1'b0;
  wire tmp265;
  assign tmp265 = (tmp262 & tmp263) | (tmp262 & tmp264) | (tmp263 & tmp264);
  wire tmp266;
  assign tmp266 = 1'b0;
  wire tmp267;
  assign tmp267 = pi5;
  wire tmp268;
  assign tmp268 = 1'b0;
  wire tmp269;
  assign tmp269 = (tmp266 & tmp267) | (tmp266 & tmp268) | (tmp267 & tmp268);
  wire tmp270;
  assign tmp270 = 1'b0;
  wire tmp271;
  assign tmp271 = 1'b0;
  wire tmp272;
  assign tmp272 = 1'b0;
  wire tmp273;
  assign tmp273 = (tmp270 & tmp271) | (tmp270 & tmp272) | (tmp271 & tmp272);
  wire tmp274;
  assign tmp274 = (tmp265 & tmp269) | (tmp265 & tmp273) | (tmp269 & tmp273);
  wire tmp275;
  assign tmp275 = 1'b0;
  wire tmp276;
  assign tmp276 = pi5;
  wire tmp277;
  assign tmp277 = 1'b0;
  wire tmp278;
  assign tmp278 = (tmp275 & tmp276) | (tmp275 & tmp277) | (tmp276 & tmp277);
  wire tmp279;
  assign tmp279 = pi5;
  wire tmp280;
  assign tmp280 = 1'b1;
  wire tmp281;
  assign tmp281 = 1'b0;
  wire tmp282;
  assign tmp282 = (tmp279 & tmp280) | (tmp279 & tmp281) | (tmp280 & tmp281);
  wire tmp283;
  assign tmp283 = 1'b0;
  wire tmp284;
  assign tmp284 = 1'b0;
  wire tmp285;
  assign tmp285 = 1'b0;
  wire tmp286;
  assign tmp286 = (tmp283 & tmp284) | (tmp283 & tmp285) | (tmp284 & tmp285);
  wire tmp287;
  assign tmp287 = (tmp278 & tmp282) | (tmp278 & tmp286) | (tmp282 & tmp286);
  wire tmp288;
  assign tmp288 = 1'b0;
  wire tmp289;
  assign tmp289 = 1'b0;
  wire tmp290;
  assign tmp290 = 1'b0;
  wire tmp291;
  assign tmp291 = (tmp288 & tmp289) | (tmp288 & tmp290) | (tmp289 & tmp290);
  wire tmp292;
  assign tmp292 = 1'b0;
  wire tmp293;
  assign tmp293 = 1'b0;
  wire tmp294;
  assign tmp294 = 1'b0;
  wire tmp295;
  assign tmp295 = (tmp292 & tmp293) | (tmp292 & tmp294) | (tmp293 & tmp294);
  wire tmp296;
  assign tmp296 = 1'b0;
  wire tmp297;
  assign tmp297 = 1'b0;
  wire tmp298;
  assign tmp298 = 1'b0;
  wire tmp299;
  assign tmp299 = (tmp296 & tmp297) | (tmp296 & tmp298) | (tmp297 & tmp298);
  wire tmp300;
  assign tmp300 = (tmp291 & tmp295) | (tmp291 & tmp299) | (tmp295 & tmp299);
  wire tmp301;
  assign tmp301 = (tmp274 & tmp287) | (tmp274 & tmp300) | (tmp287 & tmp300);
  wire tmp302;
  assign tmp302 = (tmp221 & tmp261) | (tmp221 & tmp301) | (tmp261 & tmp301);
  assign po4 = tmp302;
  wire tmp303;
  assign tmp303 = 1'b1;
  wire tmp304;
  assign tmp304 = 1'b1;
  wire tmp305;
  assign tmp305 = 1'b1;
  wire tmp306;
  assign tmp306 = (tmp303 & tmp304) | (tmp303 & tmp305) | (tmp304 & tmp305);
  wire tmp307;
  assign tmp307 = 1'b1;
  wire tmp308;
  assign tmp308 = w1;
  wire tmp309;
  assign tmp309 = pi4;
  wire tmp310;
  assign tmp310 = (tmp307 & tmp308) | (tmp307 & tmp309) | (tmp308 & tmp309);
  wire tmp311;
  assign tmp311 = 1'b1;
  wire tmp312;
  assign tmp312 = pi4;
  wire tmp313;
  assign tmp313 = pi5;
  wire tmp314;
  assign tmp314 = (tmp311 & tmp312) | (tmp311 & tmp313) | (tmp312 & tmp313);
  wire tmp315;
  assign tmp315 = (tmp306 & tmp310) | (tmp306 & tmp314) | (tmp310 & tmp314);
  wire tmp316;
  assign tmp316 = 1'b1;
  wire tmp317;
  assign tmp317 = w1;
  wire tmp318;
  assign tmp318 = pi4;
  wire tmp319;
  assign tmp319 = (tmp316 & tmp317) | (tmp316 & tmp318) | (tmp317 & tmp318);
  wire tmp320;
  assign tmp320 = w1;
  wire tmp321;
  assign tmp321 = 1'b1;
  wire tmp322;
  assign tmp322 = 1'b1;
  wire tmp323;
  assign tmp323 = (tmp320 & tmp321) | (tmp320 & tmp322) | (tmp321 & tmp322);
  wire tmp324;
  assign tmp324 = pi4;
  wire tmp325;
  assign tmp325 = 1'b1;
  wire tmp326;
  assign tmp326 = 1'b1;
  wire tmp327;
  assign tmp327 = (tmp324 & tmp325) | (tmp324 & tmp326) | (tmp325 & tmp326);
  wire tmp328;
  assign tmp328 = (tmp319 & tmp323) | (tmp319 & tmp327) | (tmp323 & tmp327);
  wire tmp329;
  assign tmp329 = 1'b1;
  wire tmp330;
  assign tmp330 = pi4;
  wire tmp331;
  assign tmp331 = pi5;
  wire tmp332;
  assign tmp332 = (tmp329 & tmp330) | (tmp329 & tmp331) | (tmp330 & tmp331);
  wire tmp333;
  assign tmp333 = pi4;
  wire tmp334;
  assign tmp334 = 1'b1;
  wire tmp335;
  assign tmp335 = 1'b1;
  wire tmp336;
  assign tmp336 = (tmp333 & tmp334) | (tmp333 & tmp335) | (tmp334 & tmp335);
  wire tmp337;
  assign tmp337 = pi5;
  wire tmp338;
  assign tmp338 = 1'b1;
  wire tmp339;
  assign tmp339 = 1'b0;
  wire tmp340;
  assign tmp340 = (tmp337 & tmp338) | (tmp337 & tmp339) | (tmp338 & tmp339);
  wire tmp341;
  assign tmp341 = (tmp332 & tmp336) | (tmp332 & tmp340) | (tmp336 & tmp340);
  wire tmp342;
  assign tmp342 = (tmp315 & tmp328) | (tmp315 & tmp341) | (tmp328 & tmp341);
  assign po5 = tmp342;
endmodule // test_each
