module test_4( pi0, pi1, pi2, pi3, pi4, po0 );
  input pi0, pi1, pi2, pi3, pi4;
  output po0;
  wire tmp0;
  assign tmp0 = 1'b1;
  wire tmp1;
  assign tmp1 = 1'b1;
  wire tmp2;
  assign tmp2 = 1'b1;
  wire tmp3;
  assign tmp3 = (tmp0 & tmp1) | (tmp0 & tmp2) | (tmp1 & tmp2);
  wire tmp4;
  assign tmp4 = 1'b1;
  wire tmp5;
  assign tmp5 = pi0;
  wire tmp6;
  assign tmp6 = pi1;
  wire tmp7;
  assign tmp7 = (tmp4 & tmp5) | (tmp4 & tmp6) | (tmp5 & tmp6);
  wire tmp8;
  assign tmp8 = 1'b1;
  wire tmp9;
  assign tmp9 = pi1;
  wire tmp10;
  assign tmp10 = pi4;
  wire tmp11;
  assign tmp11 = (tmp8 & tmp9) | (tmp8 & tmp10) | (tmp9 & tmp10);
  wire tmp12;
  assign tmp12 = (tmp3 & tmp7) | (tmp3 & tmp11) | (tmp7 & tmp11);
  wire tmp13;
  assign tmp13 = 1'b1;
  wire tmp14;
  assign tmp14 = pi0;
  wire tmp15;
  assign tmp15 = pi1;
  wire tmp16;
  assign tmp16 = (tmp13 & tmp14) | (tmp13 & tmp15) | (tmp14 & tmp15);
  wire tmp17;
  assign tmp17 = pi0;
  wire tmp18;
  assign tmp18 = 1'b1;
  wire tmp19;
  assign tmp19 = 1'b1;
  wire tmp20;
  assign tmp20 = (tmp17 & tmp18) | (tmp17 & tmp19) | (tmp18 & tmp19);
  wire tmp21;
  assign tmp21 = pi1;
  wire tmp22;
  assign tmp22 = 1'b1;
  wire tmp23;
  assign tmp23 = 1'b1;
  wire tmp24;
  assign tmp24 = (tmp21 & tmp22) | (tmp21 & tmp23) | (tmp22 & tmp23);
  wire tmp25;
  assign tmp25 = (tmp16 & tmp20) | (tmp16 & tmp24) | (tmp20 & tmp24);
  wire tmp26;
  assign tmp26 = 1'b1;
  wire tmp27;
  assign tmp27 = pi1;
  wire tmp28;
  assign tmp28 = pi4;
  wire tmp29;
  assign tmp29 = (tmp26 & tmp27) | (tmp26 & tmp28) | (tmp27 & tmp28);
  wire tmp30;
  assign tmp30 = pi1;
  wire tmp31;
  assign tmp31 = 1'b1;
  wire tmp32;
  assign tmp32 = 1'b1;
  wire tmp33;
  assign tmp33 = (tmp30 & tmp31) | (tmp30 & tmp32) | (tmp31 & tmp32);
  wire tmp34;
  assign tmp34 = pi4;
  wire tmp35;
  assign tmp35 = 1'b1;
  wire tmp36;
  assign tmp36 = 1'b0;
  wire tmp37;
  assign tmp37 = (tmp34 & tmp35) | (tmp34 & tmp36) | (tmp35 & tmp36);
  wire tmp38;
  assign tmp38 = (tmp29 & tmp33) | (tmp29 & tmp37) | (tmp33 & tmp37);
  wire tmp39;
  assign tmp39 = (tmp12 & tmp25) | (tmp12 & tmp38) | (tmp25 & tmp38);
  wire tmp40;
  assign tmp40 = 1'b1;
  wire tmp41;
  assign tmp41 = pi0;
  wire tmp42;
  assign tmp42 = pi1;
  wire tmp43;
  assign tmp43 = (tmp40 & tmp41) | (tmp40 & tmp42) | (tmp41 & tmp42);
  wire tmp44;
  assign tmp44 = pi0;
  wire tmp45;
  assign tmp45 = 1'b1;
  wire tmp46;
  assign tmp46 = 1'b1;
  wire tmp47;
  assign tmp47 = (tmp44 & tmp45) | (tmp44 & tmp46) | (tmp45 & tmp46);
  wire tmp48;
  assign tmp48 = pi1;
  wire tmp49;
  assign tmp49 = 1'b1;
  wire tmp50;
  assign tmp50 = 1'b1;
  wire tmp51;
  assign tmp51 = (tmp48 & tmp49) | (tmp48 & tmp50) | (tmp49 & tmp50);
  wire tmp52;
  assign tmp52 = (tmp43 & tmp47) | (tmp43 & tmp51) | (tmp47 & tmp51);
  wire tmp53;
  assign tmp53 = pi0;
  wire tmp54;
  assign tmp54 = 1'b1;
  wire tmp55;
  assign tmp55 = 1'b1;
  wire tmp56;
  assign tmp56 = (tmp53 & tmp54) | (tmp53 & tmp55) | (tmp54 & tmp55);
  wire tmp57;
  assign tmp57 = 1'b1;
  wire tmp58;
  assign tmp58 = 1'b1;
  wire tmp59;
  assign tmp59 = 1'b0;
  wire tmp60;
  assign tmp60 = (tmp57 & tmp58) | (tmp57 & tmp59) | (tmp58 & tmp59);
  wire tmp61;
  assign tmp61 = 1'b1;
  wire tmp62;
  assign tmp62 = 1'b0;
  wire tmp63;
  assign tmp63 = 1'b0;
  wire tmp64;
  assign tmp64 = (tmp61 & tmp62) | (tmp61 & tmp63) | (tmp62 & tmp63);
  wire tmp65;
  assign tmp65 = (tmp56 & tmp60) | (tmp56 & tmp64) | (tmp60 & tmp64);
  wire tmp66;
  assign tmp66 = pi1;
  wire tmp67;
  assign tmp67 = 1'b1;
  wire tmp68;
  assign tmp68 = 1'b1;
  wire tmp69;
  assign tmp69 = (tmp66 & tmp67) | (tmp66 & tmp68) | (tmp67 & tmp68);
  wire tmp70;
  assign tmp70 = 1'b1;
  wire tmp71;
  assign tmp71 = 1'b0;
  wire tmp72;
  assign tmp72 = 1'b0;
  wire tmp73;
  assign tmp73 = (tmp70 & tmp71) | (tmp70 & tmp72) | (tmp71 & tmp72);
  wire tmp74;
  assign tmp74 = 1'b1;
  wire tmp75;
  assign tmp75 = 1'b0;
  wire tmp76;
  assign tmp76 = 1'b0;
  wire tmp77;
  assign tmp77 = (tmp74 & tmp75) | (tmp74 & tmp76) | (tmp75 & tmp76);
  wire tmp78;
  assign tmp78 = (tmp69 & tmp73) | (tmp69 & tmp77) | (tmp73 & tmp77);
  wire tmp79;
  assign tmp79 = (tmp52 & tmp65) | (tmp52 & tmp78) | (tmp65 & tmp78);
  wire tmp80;
  assign tmp80 = 1'b1;
  wire tmp81;
  assign tmp81 = pi1;
  wire tmp82;
  assign tmp82 = pi4;
  wire tmp83;
  assign tmp83 = (tmp80 & tmp81) | (tmp80 & tmp82) | (tmp81 & tmp82);
  wire tmp84;
  assign tmp84 = pi1;
  wire tmp85;
  assign tmp85 = 1'b1;
  wire tmp86;
  assign tmp86 = 1'b1;
  wire tmp87;
  assign tmp87 = (tmp84 & tmp85) | (tmp84 & tmp86) | (tmp85 & tmp86);
  wire tmp88;
  assign tmp88 = pi4;
  wire tmp89;
  assign tmp89 = 1'b1;
  wire tmp90;
  assign tmp90 = 1'b0;
  wire tmp91;
  assign tmp91 = (tmp88 & tmp89) | (tmp88 & tmp90) | (tmp89 & tmp90);
  wire tmp92;
  assign tmp92 = (tmp83 & tmp87) | (tmp83 & tmp91) | (tmp87 & tmp91);
  wire tmp93;
  assign tmp93 = pi1;
  wire tmp94;
  assign tmp94 = 1'b1;
  wire tmp95;
  assign tmp95 = 1'b1;
  wire tmp96;
  assign tmp96 = (tmp93 & tmp94) | (tmp93 & tmp95) | (tmp94 & tmp95);
  wire tmp97;
  assign tmp97 = 1'b1;
  wire tmp98;
  assign tmp98 = 1'b0;
  wire tmp99;
  assign tmp99 = 1'b0;
  wire tmp100;
  assign tmp100 = (tmp97 & tmp98) | (tmp97 & tmp99) | (tmp98 & tmp99);
  wire tmp101;
  assign tmp101 = 1'b1;
  wire tmp102;
  assign tmp102 = 1'b0;
  wire tmp103;
  assign tmp103 = 1'b0;
  wire tmp104;
  assign tmp104 = (tmp101 & tmp102) | (tmp101 & tmp103) | (tmp102 & tmp103);
  wire tmp105;
  assign tmp105 = (tmp96 & tmp100) | (tmp96 & tmp104) | (tmp100 & tmp104);
  wire tmp106;
  assign tmp106 = pi4;
  wire tmp107;
  assign tmp107 = 1'b1;
  wire tmp108;
  assign tmp108 = 1'b0;
  wire tmp109;
  assign tmp109 = (tmp106 & tmp107) | (tmp106 & tmp108) | (tmp107 & tmp108);
  wire tmp110;
  assign tmp110 = 1'b1;
  wire tmp111;
  assign tmp111 = 1'b0;
  wire tmp112;
  assign tmp112 = 1'b0;
  wire tmp113;
  assign tmp113 = (tmp110 & tmp111) | (tmp110 & tmp112) | (tmp111 & tmp112);
  wire tmp114;
  assign tmp114 = 1'b0;
  wire tmp115;
  assign tmp115 = 1'b0;
  wire tmp116;
  assign tmp116 = 1'b0;
  wire tmp117;
  assign tmp117 = (tmp114 & tmp115) | (tmp114 & tmp116) | (tmp115 & tmp116);
  wire tmp118;
  assign tmp118 = (tmp109 & tmp113) | (tmp109 & tmp117) | (tmp113 & tmp117);
  wire tmp119;
  assign tmp119 = (tmp92 & tmp105) | (tmp92 & tmp118) | (tmp105 & tmp118);
  wire tmp120;
  assign tmp120 = (tmp39 & tmp79) | (tmp39 & tmp119) | (tmp79 & tmp119);
  wire tmp121;
  assign tmp121 = 1'b1;
  wire tmp122;
  assign tmp122 = pi0;
  wire tmp123;
  assign tmp123 = pi1;
  wire tmp124;
  assign tmp124 = (tmp121 & tmp122) | (tmp121 & tmp123) | (tmp122 & tmp123);
  wire tmp125;
  assign tmp125 = pi0;
  wire tmp126;
  assign tmp126 = 1'b1;
  wire tmp127;
  assign tmp127 = 1'b1;
  wire tmp128;
  assign tmp128 = (tmp125 & tmp126) | (tmp125 & tmp127) | (tmp126 & tmp127);
  wire tmp129;
  assign tmp129 = pi1;
  wire tmp130;
  assign tmp130 = 1'b1;
  wire tmp131;
  assign tmp131 = 1'b1;
  wire tmp132;
  assign tmp132 = (tmp129 & tmp130) | (tmp129 & tmp131) | (tmp130 & tmp131);
  wire tmp133;
  assign tmp133 = (tmp124 & tmp128) | (tmp124 & tmp132) | (tmp128 & tmp132);
  wire tmp134;
  assign tmp134 = pi0;
  wire tmp135;
  assign tmp135 = 1'b1;
  wire tmp136;
  assign tmp136 = 1'b1;
  wire tmp137;
  assign tmp137 = (tmp134 & tmp135) | (tmp134 & tmp136) | (tmp135 & tmp136);
  wire tmp138;
  assign tmp138 = 1'b1;
  wire tmp139;
  assign tmp139 = 1'b1;
  wire tmp140;
  assign tmp140 = 1'b0;
  wire tmp141;
  assign tmp141 = (tmp138 & tmp139) | (tmp138 & tmp140) | (tmp139 & tmp140);
  wire tmp142;
  assign tmp142 = 1'b1;
  wire tmp143;
  assign tmp143 = 1'b0;
  wire tmp144;
  assign tmp144 = 1'b0;
  wire tmp145;
  assign tmp145 = (tmp142 & tmp143) | (tmp142 & tmp144) | (tmp143 & tmp144);
  wire tmp146;
  assign tmp146 = (tmp137 & tmp141) | (tmp137 & tmp145) | (tmp141 & tmp145);
  wire tmp147;
  assign tmp147 = pi1;
  wire tmp148;
  assign tmp148 = 1'b1;
  wire tmp149;
  assign tmp149 = 1'b1;
  wire tmp150;
  assign tmp150 = (tmp147 & tmp148) | (tmp147 & tmp149) | (tmp148 & tmp149);
  wire tmp151;
  assign tmp151 = 1'b1;
  wire tmp152;
  assign tmp152 = 1'b0;
  wire tmp153;
  assign tmp153 = 1'b0;
  wire tmp154;
  assign tmp154 = (tmp151 & tmp152) | (tmp151 & tmp153) | (tmp152 & tmp153);
  wire tmp155;
  assign tmp155 = 1'b1;
  wire tmp156;
  assign tmp156 = 1'b0;
  wire tmp157;
  assign tmp157 = 1'b0;
  wire tmp158;
  assign tmp158 = (tmp155 & tmp156) | (tmp155 & tmp157) | (tmp156 & tmp157);
  wire tmp159;
  assign tmp159 = (tmp150 & tmp154) | (tmp150 & tmp158) | (tmp154 & tmp158);
  wire tmp160;
  assign tmp160 = (tmp133 & tmp146) | (tmp133 & tmp159) | (tmp146 & tmp159);
  wire tmp161;
  assign tmp161 = pi0;
  wire tmp162;
  assign tmp162 = 1'b1;
  wire tmp163;
  assign tmp163 = 1'b1;
  wire tmp164;
  assign tmp164 = (tmp161 & tmp162) | (tmp161 & tmp163) | (tmp162 & tmp163);
  wire tmp165;
  assign tmp165 = 1'b1;
  wire tmp166;
  assign tmp166 = 1'b1;
  wire tmp167;
  assign tmp167 = 1'b0;
  wire tmp168;
  assign tmp168 = (tmp165 & tmp166) | (tmp165 & tmp167) | (tmp166 & tmp167);
  wire tmp169;
  assign tmp169 = 1'b1;
  wire tmp170;
  assign tmp170 = 1'b0;
  wire tmp171;
  assign tmp171 = 1'b0;
  wire tmp172;
  assign tmp172 = (tmp169 & tmp170) | (tmp169 & tmp171) | (tmp170 & tmp171);
  wire tmp173;
  assign tmp173 = (tmp164 & tmp168) | (tmp164 & tmp172) | (tmp168 & tmp172);
  wire tmp174;
  assign tmp174 = 1'b1;
  wire tmp175;
  assign tmp175 = 1'b1;
  wire tmp176;
  assign tmp176 = 1'b0;
  wire tmp177;
  assign tmp177 = (tmp174 & tmp175) | (tmp174 & tmp176) | (tmp175 & tmp176);
  wire tmp178;
  assign tmp178 = 1'b1;
  wire tmp179;
  assign tmp179 = pi2;
  wire tmp180;
  assign tmp180 = pi3;
  wire tmp181;
  assign tmp181 = (tmp178 & tmp179) | (tmp178 & tmp180) | (tmp179 & tmp180);
  wire tmp182;
  assign tmp182 = 1'b0;
  wire tmp183;
  assign tmp183 = pi3;
  wire tmp184;
  assign tmp184 = 1'b0;
  wire tmp185;
  assign tmp185 = (tmp182 & tmp183) | (tmp182 & tmp184) | (tmp183 & tmp184);
  wire tmp186;
  assign tmp186 = (tmp177 & tmp181) | (tmp177 & tmp185) | (tmp181 & tmp185);
  wire tmp187;
  assign tmp187 = 1'b1;
  wire tmp188;
  assign tmp188 = 1'b0;
  wire tmp189;
  assign tmp189 = 1'b0;
  wire tmp190;
  assign tmp190 = (tmp187 & tmp188) | (tmp187 & tmp189) | (tmp188 & tmp189);
  wire tmp191;
  assign tmp191 = 1'b0;
  wire tmp192;
  assign tmp192 = pi3;
  wire tmp193;
  assign tmp193 = 1'b0;
  wire tmp194;
  assign tmp194 = (tmp191 & tmp192) | (tmp191 & tmp193) | (tmp192 & tmp193);
  wire tmp195;
  assign tmp195 = 1'b0;
  wire tmp196;
  assign tmp196 = 1'b0;
  wire tmp197;
  assign tmp197 = 1'b0;
  wire tmp198;
  assign tmp198 = (tmp195 & tmp196) | (tmp195 & tmp197) | (tmp196 & tmp197);
  wire tmp199;
  assign tmp199 = (tmp190 & tmp194) | (tmp190 & tmp198) | (tmp194 & tmp198);
  wire tmp200;
  assign tmp200 = (tmp173 & tmp186) | (tmp173 & tmp199) | (tmp186 & tmp199);
  wire tmp201;
  assign tmp201 = pi1;
  wire tmp202;
  assign tmp202 = 1'b1;
  wire tmp203;
  assign tmp203 = 1'b1;
  wire tmp204;
  assign tmp204 = (tmp201 & tmp202) | (tmp201 & tmp203) | (tmp202 & tmp203);
  wire tmp205;
  assign tmp205 = 1'b1;
  wire tmp206;
  assign tmp206 = 1'b0;
  wire tmp207;
  assign tmp207 = 1'b0;
  wire tmp208;
  assign tmp208 = (tmp205 & tmp206) | (tmp205 & tmp207) | (tmp206 & tmp207);
  wire tmp209;
  assign tmp209 = 1'b1;
  wire tmp210;
  assign tmp210 = 1'b0;
  wire tmp211;
  assign tmp211 = 1'b0;
  wire tmp212;
  assign tmp212 = (tmp209 & tmp210) | (tmp209 & tmp211) | (tmp210 & tmp211);
  wire tmp213;
  assign tmp213 = (tmp204 & tmp208) | (tmp204 & tmp212) | (tmp208 & tmp212);
  wire tmp214;
  assign tmp214 = 1'b1;
  wire tmp215;
  assign tmp215 = 1'b0;
  wire tmp216;
  assign tmp216 = 1'b0;
  wire tmp217;
  assign tmp217 = (tmp214 & tmp215) | (tmp214 & tmp216) | (tmp215 & tmp216);
  wire tmp218;
  assign tmp218 = 1'b0;
  wire tmp219;
  assign tmp219 = pi3;
  wire tmp220;
  assign tmp220 = 1'b0;
  wire tmp221;
  assign tmp221 = (tmp218 & tmp219) | (tmp218 & tmp220) | (tmp219 & tmp220);
  wire tmp222;
  assign tmp222 = 1'b0;
  wire tmp223;
  assign tmp223 = 1'b0;
  wire tmp224;
  assign tmp224 = 1'b0;
  wire tmp225;
  assign tmp225 = (tmp222 & tmp223) | (tmp222 & tmp224) | (tmp223 & tmp224);
  wire tmp226;
  assign tmp226 = (tmp217 & tmp221) | (tmp217 & tmp225) | (tmp221 & tmp225);
  wire tmp227;
  assign tmp227 = 1'b1;
  wire tmp228;
  assign tmp228 = 1'b0;
  wire tmp229;
  assign tmp229 = 1'b0;
  wire tmp230;
  assign tmp230 = (tmp227 & tmp228) | (tmp227 & tmp229) | (tmp228 & tmp229);
  wire tmp231;
  assign tmp231 = 1'b0;
  wire tmp232;
  assign tmp232 = 1'b0;
  wire tmp233;
  assign tmp233 = 1'b0;
  wire tmp234;
  assign tmp234 = (tmp231 & tmp232) | (tmp231 & tmp233) | (tmp232 & tmp233);
  wire tmp235;
  assign tmp235 = 1'b0;
  wire tmp236;
  assign tmp236 = 1'b0;
  wire tmp237;
  assign tmp237 = 1'b0;
  wire tmp238;
  assign tmp238 = (tmp235 & tmp236) | (tmp235 & tmp237) | (tmp236 & tmp237);
  wire tmp239;
  assign tmp239 = (tmp230 & tmp234) | (tmp230 & tmp238) | (tmp234 & tmp238);
  wire tmp240;
  assign tmp240 = (tmp213 & tmp226) | (tmp213 & tmp239) | (tmp226 & tmp239);
  wire tmp241;
  assign tmp241 = (tmp160 & tmp200) | (tmp160 & tmp240) | (tmp200 & tmp240);
  wire tmp242;
  assign tmp242 = 1'b1;
  wire tmp243;
  assign tmp243 = pi1;
  wire tmp244;
  assign tmp244 = pi4;
  wire tmp245;
  assign tmp245 = (tmp242 & tmp243) | (tmp242 & tmp244) | (tmp243 & tmp244);
  wire tmp246;
  assign tmp246 = pi1;
  wire tmp247;
  assign tmp247 = 1'b1;
  wire tmp248;
  assign tmp248 = 1'b1;
  wire tmp249;
  assign tmp249 = (tmp246 & tmp247) | (tmp246 & tmp248) | (tmp247 & tmp248);
  wire tmp250;
  assign tmp250 = pi4;
  wire tmp251;
  assign tmp251 = 1'b1;
  wire tmp252;
  assign tmp252 = 1'b0;
  wire tmp253;
  assign tmp253 = (tmp250 & tmp251) | (tmp250 & tmp252) | (tmp251 & tmp252);
  wire tmp254;
  assign tmp254 = (tmp245 & tmp249) | (tmp245 & tmp253) | (tmp249 & tmp253);
  wire tmp255;
  assign tmp255 = pi1;
  wire tmp256;
  assign tmp256 = 1'b1;
  wire tmp257;
  assign tmp257 = 1'b1;
  wire tmp258;
  assign tmp258 = (tmp255 & tmp256) | (tmp255 & tmp257) | (tmp256 & tmp257);
  wire tmp259;
  assign tmp259 = 1'b1;
  wire tmp260;
  assign tmp260 = 1'b0;
  wire tmp261;
  assign tmp261 = 1'b0;
  wire tmp262;
  assign tmp262 = (tmp259 & tmp260) | (tmp259 & tmp261) | (tmp260 & tmp261);
  wire tmp263;
  assign tmp263 = 1'b1;
  wire tmp264;
  assign tmp264 = 1'b0;
  wire tmp265;
  assign tmp265 = 1'b0;
  wire tmp266;
  assign tmp266 = (tmp263 & tmp264) | (tmp263 & tmp265) | (tmp264 & tmp265);
  wire tmp267;
  assign tmp267 = (tmp258 & tmp262) | (tmp258 & tmp266) | (tmp262 & tmp266);
  wire tmp268;
  assign tmp268 = pi4;
  wire tmp269;
  assign tmp269 = 1'b1;
  wire tmp270;
  assign tmp270 = 1'b0;
  wire tmp271;
  assign tmp271 = (tmp268 & tmp269) | (tmp268 & tmp270) | (tmp269 & tmp270);
  wire tmp272;
  assign tmp272 = 1'b1;
  wire tmp273;
  assign tmp273 = 1'b0;
  wire tmp274;
  assign tmp274 = 1'b0;
  wire tmp275;
  assign tmp275 = (tmp272 & tmp273) | (tmp272 & tmp274) | (tmp273 & tmp274);
  wire tmp276;
  assign tmp276 = 1'b0;
  wire tmp277;
  assign tmp277 = 1'b0;
  wire tmp278;
  assign tmp278 = 1'b0;
  wire tmp279;
  assign tmp279 = (tmp276 & tmp277) | (tmp276 & tmp278) | (tmp277 & tmp278);
  wire tmp280;
  assign tmp280 = (tmp271 & tmp275) | (tmp271 & tmp279) | (tmp275 & tmp279);
  wire tmp281;
  assign tmp281 = (tmp254 & tmp267) | (tmp254 & tmp280) | (tmp267 & tmp280);
  wire tmp282;
  assign tmp282 = pi1;
  wire tmp283;
  assign tmp283 = 1'b1;
  wire tmp284;
  assign tmp284 = 1'b1;
  wire tmp285;
  assign tmp285 = (tmp282 & tmp283) | (tmp282 & tmp284) | (tmp283 & tmp284);
  wire tmp286;
  assign tmp286 = 1'b1;
  wire tmp287;
  assign tmp287 = 1'b0;
  wire tmp288;
  assign tmp288 = 1'b0;
  wire tmp289;
  assign tmp289 = (tmp286 & tmp287) | (tmp286 & tmp288) | (tmp287 & tmp288);
  wire tmp290;
  assign tmp290 = 1'b1;
  wire tmp291;
  assign tmp291 = 1'b0;
  wire tmp292;
  assign tmp292 = 1'b0;
  wire tmp293;
  assign tmp293 = (tmp290 & tmp291) | (tmp290 & tmp292) | (tmp291 & tmp292);
  wire tmp294;
  assign tmp294 = (tmp285 & tmp289) | (tmp285 & tmp293) | (tmp289 & tmp293);
  wire tmp295;
  assign tmp295 = 1'b1;
  wire tmp296;
  assign tmp296 = 1'b0;
  wire tmp297;
  assign tmp297 = 1'b0;
  wire tmp298;
  assign tmp298 = (tmp295 & tmp296) | (tmp295 & tmp297) | (tmp296 & tmp297);
  wire tmp299;
  assign tmp299 = 1'b0;
  wire tmp300;
  assign tmp300 = pi3;
  wire tmp301;
  assign tmp301 = 1'b0;
  wire tmp302;
  assign tmp302 = (tmp299 & tmp300) | (tmp299 & tmp301) | (tmp300 & tmp301);
  wire tmp303;
  assign tmp303 = 1'b0;
  wire tmp304;
  assign tmp304 = 1'b0;
  wire tmp305;
  assign tmp305 = 1'b0;
  wire tmp306;
  assign tmp306 = (tmp303 & tmp304) | (tmp303 & tmp305) | (tmp304 & tmp305);
  wire tmp307;
  assign tmp307 = (tmp298 & tmp302) | (tmp298 & tmp306) | (tmp302 & tmp306);
  wire tmp308;
  assign tmp308 = 1'b1;
  wire tmp309;
  assign tmp309 = 1'b0;
  wire tmp310;
  assign tmp310 = 1'b0;
  wire tmp311;
  assign tmp311 = (tmp308 & tmp309) | (tmp308 & tmp310) | (tmp309 & tmp310);
  wire tmp312;
  assign tmp312 = 1'b0;
  wire tmp313;
  assign tmp313 = 1'b0;
  wire tmp314;
  assign tmp314 = 1'b0;
  wire tmp315;
  assign tmp315 = (tmp312 & tmp313) | (tmp312 & tmp314) | (tmp313 & tmp314);
  wire tmp316;
  assign tmp316 = 1'b0;
  wire tmp317;
  assign tmp317 = 1'b0;
  wire tmp318;
  assign tmp318 = 1'b0;
  wire tmp319;
  assign tmp319 = (tmp316 & tmp317) | (tmp316 & tmp318) | (tmp317 & tmp318);
  wire tmp320;
  assign tmp320 = (tmp311 & tmp315) | (tmp311 & tmp319) | (tmp315 & tmp319);
  wire tmp321;
  assign tmp321 = (tmp294 & tmp307) | (tmp294 & tmp320) | (tmp307 & tmp320);
  wire tmp322;
  assign tmp322 = pi4;
  wire tmp323;
  assign tmp323 = 1'b1;
  wire tmp324;
  assign tmp324 = 1'b0;
  wire tmp325;
  assign tmp325 = (tmp322 & tmp323) | (tmp322 & tmp324) | (tmp323 & tmp324);
  wire tmp326;
  assign tmp326 = 1'b1;
  wire tmp327;
  assign tmp327 = 1'b0;
  wire tmp328;
  assign tmp328 = 1'b0;
  wire tmp329;
  assign tmp329 = (tmp326 & tmp327) | (tmp326 & tmp328) | (tmp327 & tmp328);
  wire tmp330;
  assign tmp330 = 1'b0;
  wire tmp331;
  assign tmp331 = 1'b0;
  wire tmp332;
  assign tmp332 = 1'b0;
  wire tmp333;
  assign tmp333 = (tmp330 & tmp331) | (tmp330 & tmp332) | (tmp331 & tmp332);
  wire tmp334;
  assign tmp334 = (tmp325 & tmp329) | (tmp325 & tmp333) | (tmp329 & tmp333);
  wire tmp335;
  assign tmp335 = 1'b1;
  wire tmp336;
  assign tmp336 = 1'b0;
  wire tmp337;
  assign tmp337 = 1'b0;
  wire tmp338;
  assign tmp338 = (tmp335 & tmp336) | (tmp335 & tmp337) | (tmp336 & tmp337);
  wire tmp339;
  assign tmp339 = 1'b0;
  wire tmp340;
  assign tmp340 = 1'b0;
  wire tmp341;
  assign tmp341 = 1'b0;
  wire tmp342;
  assign tmp342 = (tmp339 & tmp340) | (tmp339 & tmp341) | (tmp340 & tmp341);
  wire tmp343;
  assign tmp343 = 1'b0;
  wire tmp344;
  assign tmp344 = 1'b0;
  wire tmp345;
  assign tmp345 = 1'b0;
  wire tmp346;
  assign tmp346 = (tmp343 & tmp344) | (tmp343 & tmp345) | (tmp344 & tmp345);
  wire tmp347;
  assign tmp347 = (tmp338 & tmp342) | (tmp338 & tmp346) | (tmp342 & tmp346);
  wire tmp348;
  assign tmp348 = 1'b0;
  wire tmp349;
  assign tmp349 = 1'b0;
  wire tmp350;
  assign tmp350 = 1'b0;
  wire tmp351;
  assign tmp351 = (tmp348 & tmp349) | (tmp348 & tmp350) | (tmp349 & tmp350);
  wire tmp352;
  assign tmp352 = 1'b0;
  wire tmp353;
  assign tmp353 = 1'b0;
  wire tmp354;
  assign tmp354 = 1'b0;
  wire tmp355;
  assign tmp355 = (tmp352 & tmp353) | (tmp352 & tmp354) | (tmp353 & tmp354);
  wire tmp356;
  assign tmp356 = 1'b0;
  wire tmp357;
  assign tmp357 = 1'b0;
  wire tmp358;
  assign tmp358 = 1'b0;
  wire tmp359;
  assign tmp359 = (tmp356 & tmp357) | (tmp356 & tmp358) | (tmp357 & tmp358);
  wire tmp360;
  assign tmp360 = (tmp351 & tmp355) | (tmp351 & tmp359) | (tmp355 & tmp359);
  wire tmp361;
  assign tmp361 = (tmp334 & tmp347) | (tmp334 & tmp360) | (tmp347 & tmp360);
  wire tmp362;
  assign tmp362 = (tmp281 & tmp321) | (tmp281 & tmp361) | (tmp321 & tmp361);
  wire tmp363;
  assign tmp363 = (tmp120 & tmp241) | (tmp120 & tmp362) | (tmp241 & tmp362);
  wire tmp364;
  assign tmp364 = 1'b1;
  wire tmp365;
  assign tmp365 = pi0;
  wire tmp366;
  assign tmp366 = pi1;
  wire tmp367;
  assign tmp367 = (tmp364 & tmp365) | (tmp364 & tmp366) | (tmp365 & tmp366);
  wire tmp368;
  assign tmp368 = pi0;
  wire tmp369;
  assign tmp369 = 1'b1;
  wire tmp370;
  assign tmp370 = 1'b1;
  wire tmp371;
  assign tmp371 = (tmp368 & tmp369) | (tmp368 & tmp370) | (tmp369 & tmp370);
  wire tmp372;
  assign tmp372 = pi1;
  wire tmp373;
  assign tmp373 = 1'b1;
  wire tmp374;
  assign tmp374 = 1'b1;
  wire tmp375;
  assign tmp375 = (tmp372 & tmp373) | (tmp372 & tmp374) | (tmp373 & tmp374);
  wire tmp376;
  assign tmp376 = (tmp367 & tmp371) | (tmp367 & tmp375) | (tmp371 & tmp375);
  wire tmp377;
  assign tmp377 = pi0;
  wire tmp378;
  assign tmp378 = 1'b1;
  wire tmp379;
  assign tmp379 = 1'b1;
  wire tmp380;
  assign tmp380 = (tmp377 & tmp378) | (tmp377 & tmp379) | (tmp378 & tmp379);
  wire tmp381;
  assign tmp381 = 1'b1;
  wire tmp382;
  assign tmp382 = 1'b1;
  wire tmp383;
  assign tmp383 = 1'b0;
  wire tmp384;
  assign tmp384 = (tmp381 & tmp382) | (tmp381 & tmp383) | (tmp382 & tmp383);
  wire tmp385;
  assign tmp385 = 1'b1;
  wire tmp386;
  assign tmp386 = 1'b0;
  wire tmp387;
  assign tmp387 = 1'b0;
  wire tmp388;
  assign tmp388 = (tmp385 & tmp386) | (tmp385 & tmp387) | (tmp386 & tmp387);
  wire tmp389;
  assign tmp389 = (tmp380 & tmp384) | (tmp380 & tmp388) | (tmp384 & tmp388);
  wire tmp390;
  assign tmp390 = pi1;
  wire tmp391;
  assign tmp391 = 1'b1;
  wire tmp392;
  assign tmp392 = 1'b1;
  wire tmp393;
  assign tmp393 = (tmp390 & tmp391) | (tmp390 & tmp392) | (tmp391 & tmp392);
  wire tmp394;
  assign tmp394 = 1'b1;
  wire tmp395;
  assign tmp395 = 1'b0;
  wire tmp396;
  assign tmp396 = 1'b0;
  wire tmp397;
  assign tmp397 = (tmp394 & tmp395) | (tmp394 & tmp396) | (tmp395 & tmp396);
  wire tmp398;
  assign tmp398 = 1'b1;
  wire tmp399;
  assign tmp399 = 1'b0;
  wire tmp400;
  assign tmp400 = 1'b0;
  wire tmp401;
  assign tmp401 = (tmp398 & tmp399) | (tmp398 & tmp400) | (tmp399 & tmp400);
  wire tmp402;
  assign tmp402 = (tmp393 & tmp397) | (tmp393 & tmp401) | (tmp397 & tmp401);
  wire tmp403;
  assign tmp403 = (tmp376 & tmp389) | (tmp376 & tmp402) | (tmp389 & tmp402);
  wire tmp404;
  assign tmp404 = pi0;
  wire tmp405;
  assign tmp405 = 1'b1;
  wire tmp406;
  assign tmp406 = 1'b1;
  wire tmp407;
  assign tmp407 = (tmp404 & tmp405) | (tmp404 & tmp406) | (tmp405 & tmp406);
  wire tmp408;
  assign tmp408 = 1'b1;
  wire tmp409;
  assign tmp409 = 1'b1;
  wire tmp410;
  assign tmp410 = 1'b0;
  wire tmp411;
  assign tmp411 = (tmp408 & tmp409) | (tmp408 & tmp410) | (tmp409 & tmp410);
  wire tmp412;
  assign tmp412 = 1'b1;
  wire tmp413;
  assign tmp413 = 1'b0;
  wire tmp414;
  assign tmp414 = 1'b0;
  wire tmp415;
  assign tmp415 = (tmp412 & tmp413) | (tmp412 & tmp414) | (tmp413 & tmp414);
  wire tmp416;
  assign tmp416 = (tmp407 & tmp411) | (tmp407 & tmp415) | (tmp411 & tmp415);
  wire tmp417;
  assign tmp417 = 1'b1;
  wire tmp418;
  assign tmp418 = 1'b1;
  wire tmp419;
  assign tmp419 = 1'b0;
  wire tmp420;
  assign tmp420 = (tmp417 & tmp418) | (tmp417 & tmp419) | (tmp418 & tmp419);
  wire tmp421;
  assign tmp421 = 1'b1;
  wire tmp422;
  assign tmp422 = pi2;
  wire tmp423;
  assign tmp423 = pi3;
  wire tmp424;
  assign tmp424 = (tmp421 & tmp422) | (tmp421 & tmp423) | (tmp422 & tmp423);
  wire tmp425;
  assign tmp425 = 1'b0;
  wire tmp426;
  assign tmp426 = pi3;
  wire tmp427;
  assign tmp427 = 1'b0;
  wire tmp428;
  assign tmp428 = (tmp425 & tmp426) | (tmp425 & tmp427) | (tmp426 & tmp427);
  wire tmp429;
  assign tmp429 = (tmp420 & tmp424) | (tmp420 & tmp428) | (tmp424 & tmp428);
  wire tmp430;
  assign tmp430 = 1'b1;
  wire tmp431;
  assign tmp431 = 1'b0;
  wire tmp432;
  assign tmp432 = 1'b0;
  wire tmp433;
  assign tmp433 = (tmp430 & tmp431) | (tmp430 & tmp432) | (tmp431 & tmp432);
  wire tmp434;
  assign tmp434 = 1'b0;
  wire tmp435;
  assign tmp435 = pi3;
  wire tmp436;
  assign tmp436 = 1'b0;
  wire tmp437;
  assign tmp437 = (tmp434 & tmp435) | (tmp434 & tmp436) | (tmp435 & tmp436);
  wire tmp438;
  assign tmp438 = 1'b0;
  wire tmp439;
  assign tmp439 = 1'b0;
  wire tmp440;
  assign tmp440 = 1'b0;
  wire tmp441;
  assign tmp441 = (tmp438 & tmp439) | (tmp438 & tmp440) | (tmp439 & tmp440);
  wire tmp442;
  assign tmp442 = (tmp433 & tmp437) | (tmp433 & tmp441) | (tmp437 & tmp441);
  wire tmp443;
  assign tmp443 = (tmp416 & tmp429) | (tmp416 & tmp442) | (tmp429 & tmp442);
  wire tmp444;
  assign tmp444 = pi1;
  wire tmp445;
  assign tmp445 = 1'b1;
  wire tmp446;
  assign tmp446 = 1'b1;
  wire tmp447;
  assign tmp447 = (tmp444 & tmp445) | (tmp444 & tmp446) | (tmp445 & tmp446);
  wire tmp448;
  assign tmp448 = 1'b1;
  wire tmp449;
  assign tmp449 = 1'b0;
  wire tmp450;
  assign tmp450 = 1'b0;
  wire tmp451;
  assign tmp451 = (tmp448 & tmp449) | (tmp448 & tmp450) | (tmp449 & tmp450);
  wire tmp452;
  assign tmp452 = 1'b1;
  wire tmp453;
  assign tmp453 = 1'b0;
  wire tmp454;
  assign tmp454 = 1'b0;
  wire tmp455;
  assign tmp455 = (tmp452 & tmp453) | (tmp452 & tmp454) | (tmp453 & tmp454);
  wire tmp456;
  assign tmp456 = (tmp447 & tmp451) | (tmp447 & tmp455) | (tmp451 & tmp455);
  wire tmp457;
  assign tmp457 = 1'b1;
  wire tmp458;
  assign tmp458 = 1'b0;
  wire tmp459;
  assign tmp459 = 1'b0;
  wire tmp460;
  assign tmp460 = (tmp457 & tmp458) | (tmp457 & tmp459) | (tmp458 & tmp459);
  wire tmp461;
  assign tmp461 = 1'b0;
  wire tmp462;
  assign tmp462 = pi3;
  wire tmp463;
  assign tmp463 = 1'b0;
  wire tmp464;
  assign tmp464 = (tmp461 & tmp462) | (tmp461 & tmp463) | (tmp462 & tmp463);
  wire tmp465;
  assign tmp465 = 1'b0;
  wire tmp466;
  assign tmp466 = 1'b0;
  wire tmp467;
  assign tmp467 = 1'b0;
  wire tmp468;
  assign tmp468 = (tmp465 & tmp466) | (tmp465 & tmp467) | (tmp466 & tmp467);
  wire tmp469;
  assign tmp469 = (tmp460 & tmp464) | (tmp460 & tmp468) | (tmp464 & tmp468);
  wire tmp470;
  assign tmp470 = 1'b1;
  wire tmp471;
  assign tmp471 = 1'b0;
  wire tmp472;
  assign tmp472 = 1'b0;
  wire tmp473;
  assign tmp473 = (tmp470 & tmp471) | (tmp470 & tmp472) | (tmp471 & tmp472);
  wire tmp474;
  assign tmp474 = 1'b0;
  wire tmp475;
  assign tmp475 = 1'b0;
  wire tmp476;
  assign tmp476 = 1'b0;
  wire tmp477;
  assign tmp477 = (tmp474 & tmp475) | (tmp474 & tmp476) | (tmp475 & tmp476);
  wire tmp478;
  assign tmp478 = 1'b0;
  wire tmp479;
  assign tmp479 = 1'b0;
  wire tmp480;
  assign tmp480 = 1'b0;
  wire tmp481;
  assign tmp481 = (tmp478 & tmp479) | (tmp478 & tmp480) | (tmp479 & tmp480);
  wire tmp482;
  assign tmp482 = (tmp473 & tmp477) | (tmp473 & tmp481) | (tmp477 & tmp481);
  wire tmp483;
  assign tmp483 = (tmp456 & tmp469) | (tmp456 & tmp482) | (tmp469 & tmp482);
  wire tmp484;
  assign tmp484 = (tmp403 & tmp443) | (tmp403 & tmp483) | (tmp443 & tmp483);
  wire tmp485;
  assign tmp485 = pi0;
  wire tmp486;
  assign tmp486 = 1'b1;
  wire tmp487;
  assign tmp487 = 1'b1;
  wire tmp488;
  assign tmp488 = (tmp485 & tmp486) | (tmp485 & tmp487) | (tmp486 & tmp487);
  wire tmp489;
  assign tmp489 = 1'b1;
  wire tmp490;
  assign tmp490 = 1'b1;
  wire tmp491;
  assign tmp491 = 1'b0;
  wire tmp492;
  assign tmp492 = (tmp489 & tmp490) | (tmp489 & tmp491) | (tmp490 & tmp491);
  wire tmp493;
  assign tmp493 = 1'b1;
  wire tmp494;
  assign tmp494 = 1'b0;
  wire tmp495;
  assign tmp495 = 1'b0;
  wire tmp496;
  assign tmp496 = (tmp493 & tmp494) | (tmp493 & tmp495) | (tmp494 & tmp495);
  wire tmp497;
  assign tmp497 = (tmp488 & tmp492) | (tmp488 & tmp496) | (tmp492 & tmp496);
  wire tmp498;
  assign tmp498 = 1'b1;
  wire tmp499;
  assign tmp499 = 1'b1;
  wire tmp500;
  assign tmp500 = 1'b0;
  wire tmp501;
  assign tmp501 = (tmp498 & tmp499) | (tmp498 & tmp500) | (tmp499 & tmp500);
  wire tmp502;
  assign tmp502 = 1'b1;
  wire tmp503;
  assign tmp503 = pi2;
  wire tmp504;
  assign tmp504 = pi3;
  wire tmp505;
  assign tmp505 = (tmp502 & tmp503) | (tmp502 & tmp504) | (tmp503 & tmp504);
  wire tmp506;
  assign tmp506 = 1'b0;
  wire tmp507;
  assign tmp507 = pi3;
  wire tmp508;
  assign tmp508 = 1'b0;
  wire tmp509;
  assign tmp509 = (tmp506 & tmp507) | (tmp506 & tmp508) | (tmp507 & tmp508);
  wire tmp510;
  assign tmp510 = (tmp501 & tmp505) | (tmp501 & tmp509) | (tmp505 & tmp509);
  wire tmp511;
  assign tmp511 = 1'b1;
  wire tmp512;
  assign tmp512 = 1'b0;
  wire tmp513;
  assign tmp513 = 1'b0;
  wire tmp514;
  assign tmp514 = (tmp511 & tmp512) | (tmp511 & tmp513) | (tmp512 & tmp513);
  wire tmp515;
  assign tmp515 = 1'b0;
  wire tmp516;
  assign tmp516 = pi3;
  wire tmp517;
  assign tmp517 = 1'b0;
  wire tmp518;
  assign tmp518 = (tmp515 & tmp516) | (tmp515 & tmp517) | (tmp516 & tmp517);
  wire tmp519;
  assign tmp519 = 1'b0;
  wire tmp520;
  assign tmp520 = 1'b0;
  wire tmp521;
  assign tmp521 = 1'b0;
  wire tmp522;
  assign tmp522 = (tmp519 & tmp520) | (tmp519 & tmp521) | (tmp520 & tmp521);
  wire tmp523;
  assign tmp523 = (tmp514 & tmp518) | (tmp514 & tmp522) | (tmp518 & tmp522);
  wire tmp524;
  assign tmp524 = (tmp497 & tmp510) | (tmp497 & tmp523) | (tmp510 & tmp523);
  wire tmp525;
  assign tmp525 = 1'b1;
  wire tmp526;
  assign tmp526 = 1'b1;
  wire tmp527;
  assign tmp527 = 1'b0;
  wire tmp528;
  assign tmp528 = (tmp525 & tmp526) | (tmp525 & tmp527) | (tmp526 & tmp527);
  wire tmp529;
  assign tmp529 = 1'b1;
  wire tmp530;
  assign tmp530 = pi2;
  wire tmp531;
  assign tmp531 = pi3;
  wire tmp532;
  assign tmp532 = (tmp529 & tmp530) | (tmp529 & tmp531) | (tmp530 & tmp531);
  wire tmp533;
  assign tmp533 = 1'b0;
  wire tmp534;
  assign tmp534 = pi3;
  wire tmp535;
  assign tmp535 = 1'b0;
  wire tmp536;
  assign tmp536 = (tmp533 & tmp534) | (tmp533 & tmp535) | (tmp534 & tmp535);
  wire tmp537;
  assign tmp537 = (tmp528 & tmp532) | (tmp528 & tmp536) | (tmp532 & tmp536);
  wire tmp538;
  assign tmp538 = 1'b1;
  wire tmp539;
  assign tmp539 = pi2;
  wire tmp540;
  assign tmp540 = pi3;
  wire tmp541;
  assign tmp541 = (tmp538 & tmp539) | (tmp538 & tmp540) | (tmp539 & tmp540);
  wire tmp542;
  assign tmp542 = pi2;
  wire tmp543;
  assign tmp543 = 1'b1;
  wire tmp544;
  assign tmp544 = 1'b1;
  wire tmp545;
  assign tmp545 = (tmp542 & tmp543) | (tmp542 & tmp544) | (tmp543 & tmp544);
  wire tmp546;
  assign tmp546 = pi3;
  wire tmp547;
  assign tmp547 = 1'b1;
  wire tmp548;
  assign tmp548 = 1'b0;
  wire tmp549;
  assign tmp549 = (tmp546 & tmp547) | (tmp546 & tmp548) | (tmp547 & tmp548);
  wire tmp550;
  assign tmp550 = (tmp541 & tmp545) | (tmp541 & tmp549) | (tmp545 & tmp549);
  wire tmp551;
  assign tmp551 = 1'b0;
  wire tmp552;
  assign tmp552 = pi3;
  wire tmp553;
  assign tmp553 = 1'b0;
  wire tmp554;
  assign tmp554 = (tmp551 & tmp552) | (tmp551 & tmp553) | (tmp552 & tmp553);
  wire tmp555;
  assign tmp555 = pi3;
  wire tmp556;
  assign tmp556 = 1'b1;
  wire tmp557;
  assign tmp557 = 1'b0;
  wire tmp558;
  assign tmp558 = (tmp555 & tmp556) | (tmp555 & tmp557) | (tmp556 & tmp557);
  wire tmp559;
  assign tmp559 = 1'b0;
  wire tmp560;
  assign tmp560 = 1'b0;
  wire tmp561;
  assign tmp561 = 1'b0;
  wire tmp562;
  assign tmp562 = (tmp559 & tmp560) | (tmp559 & tmp561) | (tmp560 & tmp561);
  wire tmp563;
  assign tmp563 = (tmp554 & tmp558) | (tmp554 & tmp562) | (tmp558 & tmp562);
  wire tmp564;
  assign tmp564 = (tmp537 & tmp550) | (tmp537 & tmp563) | (tmp550 & tmp563);
  wire tmp565;
  assign tmp565 = 1'b1;
  wire tmp566;
  assign tmp566 = 1'b0;
  wire tmp567;
  assign tmp567 = 1'b0;
  wire tmp568;
  assign tmp568 = (tmp565 & tmp566) | (tmp565 & tmp567) | (tmp566 & tmp567);
  wire tmp569;
  assign tmp569 = 1'b0;
  wire tmp570;
  assign tmp570 = pi3;
  wire tmp571;
  assign tmp571 = 1'b0;
  wire tmp572;
  assign tmp572 = (tmp569 & tmp570) | (tmp569 & tmp571) | (tmp570 & tmp571);
  wire tmp573;
  assign tmp573 = 1'b0;
  wire tmp574;
  assign tmp574 = 1'b0;
  wire tmp575;
  assign tmp575 = 1'b0;
  wire tmp576;
  assign tmp576 = (tmp573 & tmp574) | (tmp573 & tmp575) | (tmp574 & tmp575);
  wire tmp577;
  assign tmp577 = (tmp568 & tmp572) | (tmp568 & tmp576) | (tmp572 & tmp576);
  wire tmp578;
  assign tmp578 = 1'b0;
  wire tmp579;
  assign tmp579 = pi3;
  wire tmp580;
  assign tmp580 = 1'b0;
  wire tmp581;
  assign tmp581 = (tmp578 & tmp579) | (tmp578 & tmp580) | (tmp579 & tmp580);
  wire tmp582;
  assign tmp582 = pi3;
  wire tmp583;
  assign tmp583 = 1'b1;
  wire tmp584;
  assign tmp584 = 1'b0;
  wire tmp585;
  assign tmp585 = (tmp582 & tmp583) | (tmp582 & tmp584) | (tmp583 & tmp584);
  wire tmp586;
  assign tmp586 = 1'b0;
  wire tmp587;
  assign tmp587 = 1'b0;
  wire tmp588;
  assign tmp588 = 1'b0;
  wire tmp589;
  assign tmp589 = (tmp586 & tmp587) | (tmp586 & tmp588) | (tmp587 & tmp588);
  wire tmp590;
  assign tmp590 = (tmp581 & tmp585) | (tmp581 & tmp589) | (tmp585 & tmp589);
  wire tmp591;
  assign tmp591 = 1'b0;
  wire tmp592;
  assign tmp592 = 1'b0;
  wire tmp593;
  assign tmp593 = 1'b0;
  wire tmp594;
  assign tmp594 = (tmp591 & tmp592) | (tmp591 & tmp593) | (tmp592 & tmp593);
  wire tmp595;
  assign tmp595 = 1'b0;
  wire tmp596;
  assign tmp596 = 1'b0;
  wire tmp597;
  assign tmp597 = 1'b0;
  wire tmp598;
  assign tmp598 = (tmp595 & tmp596) | (tmp595 & tmp597) | (tmp596 & tmp597);
  wire tmp599;
  assign tmp599 = 1'b0;
  wire tmp600;
  assign tmp600 = 1'b0;
  wire tmp601;
  assign tmp601 = 1'b0;
  wire tmp602;
  assign tmp602 = (tmp599 & tmp600) | (tmp599 & tmp601) | (tmp600 & tmp601);
  wire tmp603;
  assign tmp603 = (tmp594 & tmp598) | (tmp594 & tmp602) | (tmp598 & tmp602);
  wire tmp604;
  assign tmp604 = (tmp577 & tmp590) | (tmp577 & tmp603) | (tmp590 & tmp603);
  wire tmp605;
  assign tmp605 = (tmp524 & tmp564) | (tmp524 & tmp604) | (tmp564 & tmp604);
  wire tmp606;
  assign tmp606 = pi1;
  wire tmp607;
  assign tmp607 = 1'b1;
  wire tmp608;
  assign tmp608 = 1'b1;
  wire tmp609;
  assign tmp609 = (tmp606 & tmp607) | (tmp606 & tmp608) | (tmp607 & tmp608);
  wire tmp610;
  assign tmp610 = 1'b1;
  wire tmp611;
  assign tmp611 = 1'b0;
  wire tmp612;
  assign tmp612 = 1'b0;
  wire tmp613;
  assign tmp613 = (tmp610 & tmp611) | (tmp610 & tmp612) | (tmp611 & tmp612);
  wire tmp614;
  assign tmp614 = 1'b1;
  wire tmp615;
  assign tmp615 = 1'b0;
  wire tmp616;
  assign tmp616 = 1'b0;
  wire tmp617;
  assign tmp617 = (tmp614 & tmp615) | (tmp614 & tmp616) | (tmp615 & tmp616);
  wire tmp618;
  assign tmp618 = (tmp609 & tmp613) | (tmp609 & tmp617) | (tmp613 & tmp617);
  wire tmp619;
  assign tmp619 = 1'b1;
  wire tmp620;
  assign tmp620 = 1'b0;
  wire tmp621;
  assign tmp621 = 1'b0;
  wire tmp622;
  assign tmp622 = (tmp619 & tmp620) | (tmp619 & tmp621) | (tmp620 & tmp621);
  wire tmp623;
  assign tmp623 = 1'b0;
  wire tmp624;
  assign tmp624 = pi3;
  wire tmp625;
  assign tmp625 = 1'b0;
  wire tmp626;
  assign tmp626 = (tmp623 & tmp624) | (tmp623 & tmp625) | (tmp624 & tmp625);
  wire tmp627;
  assign tmp627 = 1'b0;
  wire tmp628;
  assign tmp628 = 1'b0;
  wire tmp629;
  assign tmp629 = 1'b0;
  wire tmp630;
  assign tmp630 = (tmp627 & tmp628) | (tmp627 & tmp629) | (tmp628 & tmp629);
  wire tmp631;
  assign tmp631 = (tmp622 & tmp626) | (tmp622 & tmp630) | (tmp626 & tmp630);
  wire tmp632;
  assign tmp632 = 1'b1;
  wire tmp633;
  assign tmp633 = 1'b0;
  wire tmp634;
  assign tmp634 = 1'b0;
  wire tmp635;
  assign tmp635 = (tmp632 & tmp633) | (tmp632 & tmp634) | (tmp633 & tmp634);
  wire tmp636;
  assign tmp636 = 1'b0;
  wire tmp637;
  assign tmp637 = 1'b0;
  wire tmp638;
  assign tmp638 = 1'b0;
  wire tmp639;
  assign tmp639 = (tmp636 & tmp637) | (tmp636 & tmp638) | (tmp637 & tmp638);
  wire tmp640;
  assign tmp640 = 1'b0;
  wire tmp641;
  assign tmp641 = 1'b0;
  wire tmp642;
  assign tmp642 = 1'b0;
  wire tmp643;
  assign tmp643 = (tmp640 & tmp641) | (tmp640 & tmp642) | (tmp641 & tmp642);
  wire tmp644;
  assign tmp644 = (tmp635 & tmp639) | (tmp635 & tmp643) | (tmp639 & tmp643);
  wire tmp645;
  assign tmp645 = (tmp618 & tmp631) | (tmp618 & tmp644) | (tmp631 & tmp644);
  wire tmp646;
  assign tmp646 = 1'b1;
  wire tmp647;
  assign tmp647 = 1'b0;
  wire tmp648;
  assign tmp648 = 1'b0;
  wire tmp649;
  assign tmp649 = (tmp646 & tmp647) | (tmp646 & tmp648) | (tmp647 & tmp648);
  wire tmp650;
  assign tmp650 = 1'b0;
  wire tmp651;
  assign tmp651 = pi3;
  wire tmp652;
  assign tmp652 = 1'b0;
  wire tmp653;
  assign tmp653 = (tmp650 & tmp651) | (tmp650 & tmp652) | (tmp651 & tmp652);
  wire tmp654;
  assign tmp654 = 1'b0;
  wire tmp655;
  assign tmp655 = 1'b0;
  wire tmp656;
  assign tmp656 = 1'b0;
  wire tmp657;
  assign tmp657 = (tmp654 & tmp655) | (tmp654 & tmp656) | (tmp655 & tmp656);
  wire tmp658;
  assign tmp658 = (tmp649 & tmp653) | (tmp649 & tmp657) | (tmp653 & tmp657);
  wire tmp659;
  assign tmp659 = 1'b0;
  wire tmp660;
  assign tmp660 = pi3;
  wire tmp661;
  assign tmp661 = 1'b0;
  wire tmp662;
  assign tmp662 = (tmp659 & tmp660) | (tmp659 & tmp661) | (tmp660 & tmp661);
  wire tmp663;
  assign tmp663 = pi3;
  wire tmp664;
  assign tmp664 = 1'b1;
  wire tmp665;
  assign tmp665 = 1'b0;
  wire tmp666;
  assign tmp666 = (tmp663 & tmp664) | (tmp663 & tmp665) | (tmp664 & tmp665);
  wire tmp667;
  assign tmp667 = 1'b0;
  wire tmp668;
  assign tmp668 = 1'b0;
  wire tmp669;
  assign tmp669 = 1'b0;
  wire tmp670;
  assign tmp670 = (tmp667 & tmp668) | (tmp667 & tmp669) | (tmp668 & tmp669);
  wire tmp671;
  assign tmp671 = (tmp662 & tmp666) | (tmp662 & tmp670) | (tmp666 & tmp670);
  wire tmp672;
  assign tmp672 = 1'b0;
  wire tmp673;
  assign tmp673 = 1'b0;
  wire tmp674;
  assign tmp674 = 1'b0;
  wire tmp675;
  assign tmp675 = (tmp672 & tmp673) | (tmp672 & tmp674) | (tmp673 & tmp674);
  wire tmp676;
  assign tmp676 = 1'b0;
  wire tmp677;
  assign tmp677 = 1'b0;
  wire tmp678;
  assign tmp678 = 1'b0;
  wire tmp679;
  assign tmp679 = (tmp676 & tmp677) | (tmp676 & tmp678) | (tmp677 & tmp678);
  wire tmp680;
  assign tmp680 = 1'b0;
  wire tmp681;
  assign tmp681 = 1'b0;
  wire tmp682;
  assign tmp682 = 1'b0;
  wire tmp683;
  assign tmp683 = (tmp680 & tmp681) | (tmp680 & tmp682) | (tmp681 & tmp682);
  wire tmp684;
  assign tmp684 = (tmp675 & tmp679) | (tmp675 & tmp683) | (tmp679 & tmp683);
  wire tmp685;
  assign tmp685 = (tmp658 & tmp671) | (tmp658 & tmp684) | (tmp671 & tmp684);
  wire tmp686;
  assign tmp686 = 1'b1;
  wire tmp687;
  assign tmp687 = 1'b0;
  wire tmp688;
  assign tmp688 = 1'b0;
  wire tmp689;
  assign tmp689 = (tmp686 & tmp687) | (tmp686 & tmp688) | (tmp687 & tmp688);
  wire tmp690;
  assign tmp690 = 1'b0;
  wire tmp691;
  assign tmp691 = 1'b0;
  wire tmp692;
  assign tmp692 = 1'b0;
  wire tmp693;
  assign tmp693 = (tmp690 & tmp691) | (tmp690 & tmp692) | (tmp691 & tmp692);
  wire tmp694;
  assign tmp694 = 1'b0;
  wire tmp695;
  assign tmp695 = 1'b0;
  wire tmp696;
  assign tmp696 = 1'b0;
  wire tmp697;
  assign tmp697 = (tmp694 & tmp695) | (tmp694 & tmp696) | (tmp695 & tmp696);
  wire tmp698;
  assign tmp698 = (tmp689 & tmp693) | (tmp689 & tmp697) | (tmp693 & tmp697);
  wire tmp699;
  assign tmp699 = 1'b0;
  wire tmp700;
  assign tmp700 = 1'b0;
  wire tmp701;
  assign tmp701 = 1'b0;
  wire tmp702;
  assign tmp702 = (tmp699 & tmp700) | (tmp699 & tmp701) | (tmp700 & tmp701);
  wire tmp703;
  assign tmp703 = 1'b0;
  wire tmp704;
  assign tmp704 = 1'b0;
  wire tmp705;
  assign tmp705 = 1'b0;
  wire tmp706;
  assign tmp706 = (tmp703 & tmp704) | (tmp703 & tmp705) | (tmp704 & tmp705);
  wire tmp707;
  assign tmp707 = 1'b0;
  wire tmp708;
  assign tmp708 = 1'b0;
  wire tmp709;
  assign tmp709 = 1'b0;
  wire tmp710;
  assign tmp710 = (tmp707 & tmp708) | (tmp707 & tmp709) | (tmp708 & tmp709);
  wire tmp711;
  assign tmp711 = (tmp702 & tmp706) | (tmp702 & tmp710) | (tmp706 & tmp710);
  wire tmp712;
  assign tmp712 = 1'b0;
  wire tmp713;
  assign tmp713 = 1'b0;
  wire tmp714;
  assign tmp714 = 1'b0;
  wire tmp715;
  assign tmp715 = (tmp712 & tmp713) | (tmp712 & tmp714) | (tmp713 & tmp714);
  wire tmp716;
  assign tmp716 = 1'b0;
  wire tmp717;
  assign tmp717 = 1'b0;
  wire tmp718;
  assign tmp718 = 1'b0;
  wire tmp719;
  assign tmp719 = (tmp716 & tmp717) | (tmp716 & tmp718) | (tmp717 & tmp718);
  wire tmp720;
  assign tmp720 = 1'b0;
  wire tmp721;
  assign tmp721 = 1'b0;
  wire tmp722;
  assign tmp722 = 1'b0;
  wire tmp723;
  assign tmp723 = (tmp720 & tmp721) | (tmp720 & tmp722) | (tmp721 & tmp722);
  wire tmp724;
  assign tmp724 = (tmp715 & tmp719) | (tmp715 & tmp723) | (tmp719 & tmp723);
  wire tmp725;
  assign tmp725 = (tmp698 & tmp711) | (tmp698 & tmp724) | (tmp711 & tmp724);
  wire tmp726;
  assign tmp726 = (tmp645 & tmp685) | (tmp645 & tmp725) | (tmp685 & tmp725);
  wire tmp727;
  assign tmp727 = (tmp484 & tmp605) | (tmp484 & tmp726) | (tmp605 & tmp726);
  wire tmp728;
  assign tmp728 = 1'b1;
  wire tmp729;
  assign tmp729 = pi1;
  wire tmp730;
  assign tmp730 = pi4;
  wire tmp731;
  assign tmp731 = (tmp728 & tmp729) | (tmp728 & tmp730) | (tmp729 & tmp730);
  wire tmp732;
  assign tmp732 = pi1;
  wire tmp733;
  assign tmp733 = 1'b1;
  wire tmp734;
  assign tmp734 = 1'b1;
  wire tmp735;
  assign tmp735 = (tmp732 & tmp733) | (tmp732 & tmp734) | (tmp733 & tmp734);
  wire tmp736;
  assign tmp736 = pi4;
  wire tmp737;
  assign tmp737 = 1'b1;
  wire tmp738;
  assign tmp738 = 1'b0;
  wire tmp739;
  assign tmp739 = (tmp736 & tmp737) | (tmp736 & tmp738) | (tmp737 & tmp738);
  wire tmp740;
  assign tmp740 = (tmp731 & tmp735) | (tmp731 & tmp739) | (tmp735 & tmp739);
  wire tmp741;
  assign tmp741 = pi1;
  wire tmp742;
  assign tmp742 = 1'b1;
  wire tmp743;
  assign tmp743 = 1'b1;
  wire tmp744;
  assign tmp744 = (tmp741 & tmp742) | (tmp741 & tmp743) | (tmp742 & tmp743);
  wire tmp745;
  assign tmp745 = 1'b1;
  wire tmp746;
  assign tmp746 = 1'b0;
  wire tmp747;
  assign tmp747 = 1'b0;
  wire tmp748;
  assign tmp748 = (tmp745 & tmp746) | (tmp745 & tmp747) | (tmp746 & tmp747);
  wire tmp749;
  assign tmp749 = 1'b1;
  wire tmp750;
  assign tmp750 = 1'b0;
  wire tmp751;
  assign tmp751 = 1'b0;
  wire tmp752;
  assign tmp752 = (tmp749 & tmp750) | (tmp749 & tmp751) | (tmp750 & tmp751);
  wire tmp753;
  assign tmp753 = (tmp744 & tmp748) | (tmp744 & tmp752) | (tmp748 & tmp752);
  wire tmp754;
  assign tmp754 = pi4;
  wire tmp755;
  assign tmp755 = 1'b1;
  wire tmp756;
  assign tmp756 = 1'b0;
  wire tmp757;
  assign tmp757 = (tmp754 & tmp755) | (tmp754 & tmp756) | (tmp755 & tmp756);
  wire tmp758;
  assign tmp758 = 1'b1;
  wire tmp759;
  assign tmp759 = 1'b0;
  wire tmp760;
  assign tmp760 = 1'b0;
  wire tmp761;
  assign tmp761 = (tmp758 & tmp759) | (tmp758 & tmp760) | (tmp759 & tmp760);
  wire tmp762;
  assign tmp762 = 1'b0;
  wire tmp763;
  assign tmp763 = 1'b0;
  wire tmp764;
  assign tmp764 = 1'b0;
  wire tmp765;
  assign tmp765 = (tmp762 & tmp763) | (tmp762 & tmp764) | (tmp763 & tmp764);
  wire tmp766;
  assign tmp766 = (tmp757 & tmp761) | (tmp757 & tmp765) | (tmp761 & tmp765);
  wire tmp767;
  assign tmp767 = (tmp740 & tmp753) | (tmp740 & tmp766) | (tmp753 & tmp766);
  wire tmp768;
  assign tmp768 = pi1;
  wire tmp769;
  assign tmp769 = 1'b1;
  wire tmp770;
  assign tmp770 = 1'b1;
  wire tmp771;
  assign tmp771 = (tmp768 & tmp769) | (tmp768 & tmp770) | (tmp769 & tmp770);
  wire tmp772;
  assign tmp772 = 1'b1;
  wire tmp773;
  assign tmp773 = 1'b0;
  wire tmp774;
  assign tmp774 = 1'b0;
  wire tmp775;
  assign tmp775 = (tmp772 & tmp773) | (tmp772 & tmp774) | (tmp773 & tmp774);
  wire tmp776;
  assign tmp776 = 1'b1;
  wire tmp777;
  assign tmp777 = 1'b0;
  wire tmp778;
  assign tmp778 = 1'b0;
  wire tmp779;
  assign tmp779 = (tmp776 & tmp777) | (tmp776 & tmp778) | (tmp777 & tmp778);
  wire tmp780;
  assign tmp780 = (tmp771 & tmp775) | (tmp771 & tmp779) | (tmp775 & tmp779);
  wire tmp781;
  assign tmp781 = 1'b1;
  wire tmp782;
  assign tmp782 = 1'b0;
  wire tmp783;
  assign tmp783 = 1'b0;
  wire tmp784;
  assign tmp784 = (tmp781 & tmp782) | (tmp781 & tmp783) | (tmp782 & tmp783);
  wire tmp785;
  assign tmp785 = 1'b0;
  wire tmp786;
  assign tmp786 = pi3;
  wire tmp787;
  assign tmp787 = 1'b0;
  wire tmp788;
  assign tmp788 = (tmp785 & tmp786) | (tmp785 & tmp787) | (tmp786 & tmp787);
  wire tmp789;
  assign tmp789 = 1'b0;
  wire tmp790;
  assign tmp790 = 1'b0;
  wire tmp791;
  assign tmp791 = 1'b0;
  wire tmp792;
  assign tmp792 = (tmp789 & tmp790) | (tmp789 & tmp791) | (tmp790 & tmp791);
  wire tmp793;
  assign tmp793 = (tmp784 & tmp788) | (tmp784 & tmp792) | (tmp788 & tmp792);
  wire tmp794;
  assign tmp794 = 1'b1;
  wire tmp795;
  assign tmp795 = 1'b0;
  wire tmp796;
  assign tmp796 = 1'b0;
  wire tmp797;
  assign tmp797 = (tmp794 & tmp795) | (tmp794 & tmp796) | (tmp795 & tmp796);
  wire tmp798;
  assign tmp798 = 1'b0;
  wire tmp799;
  assign tmp799 = 1'b0;
  wire tmp800;
  assign tmp800 = 1'b0;
  wire tmp801;
  assign tmp801 = (tmp798 & tmp799) | (tmp798 & tmp800) | (tmp799 & tmp800);
  wire tmp802;
  assign tmp802 = 1'b0;
  wire tmp803;
  assign tmp803 = 1'b0;
  wire tmp804;
  assign tmp804 = 1'b0;
  wire tmp805;
  assign tmp805 = (tmp802 & tmp803) | (tmp802 & tmp804) | (tmp803 & tmp804);
  wire tmp806;
  assign tmp806 = (tmp797 & tmp801) | (tmp797 & tmp805) | (tmp801 & tmp805);
  wire tmp807;
  assign tmp807 = (tmp780 & tmp793) | (tmp780 & tmp806) | (tmp793 & tmp806);
  wire tmp808;
  assign tmp808 = pi4;
  wire tmp809;
  assign tmp809 = 1'b1;
  wire tmp810;
  assign tmp810 = 1'b0;
  wire tmp811;
  assign tmp811 = (tmp808 & tmp809) | (tmp808 & tmp810) | (tmp809 & tmp810);
  wire tmp812;
  assign tmp812 = 1'b1;
  wire tmp813;
  assign tmp813 = 1'b0;
  wire tmp814;
  assign tmp814 = 1'b0;
  wire tmp815;
  assign tmp815 = (tmp812 & tmp813) | (tmp812 & tmp814) | (tmp813 & tmp814);
  wire tmp816;
  assign tmp816 = 1'b0;
  wire tmp817;
  assign tmp817 = 1'b0;
  wire tmp818;
  assign tmp818 = 1'b0;
  wire tmp819;
  assign tmp819 = (tmp816 & tmp817) | (tmp816 & tmp818) | (tmp817 & tmp818);
  wire tmp820;
  assign tmp820 = (tmp811 & tmp815) | (tmp811 & tmp819) | (tmp815 & tmp819);
  wire tmp821;
  assign tmp821 = 1'b1;
  wire tmp822;
  assign tmp822 = 1'b0;
  wire tmp823;
  assign tmp823 = 1'b0;
  wire tmp824;
  assign tmp824 = (tmp821 & tmp822) | (tmp821 & tmp823) | (tmp822 & tmp823);
  wire tmp825;
  assign tmp825 = 1'b0;
  wire tmp826;
  assign tmp826 = 1'b0;
  wire tmp827;
  assign tmp827 = 1'b0;
  wire tmp828;
  assign tmp828 = (tmp825 & tmp826) | (tmp825 & tmp827) | (tmp826 & tmp827);
  wire tmp829;
  assign tmp829 = 1'b0;
  wire tmp830;
  assign tmp830 = 1'b0;
  wire tmp831;
  assign tmp831 = 1'b0;
  wire tmp832;
  assign tmp832 = (tmp829 & tmp830) | (tmp829 & tmp831) | (tmp830 & tmp831);
  wire tmp833;
  assign tmp833 = (tmp824 & tmp828) | (tmp824 & tmp832) | (tmp828 & tmp832);
  wire tmp834;
  assign tmp834 = 1'b0;
  wire tmp835;
  assign tmp835 = 1'b0;
  wire tmp836;
  assign tmp836 = 1'b0;
  wire tmp837;
  assign tmp837 = (tmp834 & tmp835) | (tmp834 & tmp836) | (tmp835 & tmp836);
  wire tmp838;
  assign tmp838 = 1'b0;
  wire tmp839;
  assign tmp839 = 1'b0;
  wire tmp840;
  assign tmp840 = 1'b0;
  wire tmp841;
  assign tmp841 = (tmp838 & tmp839) | (tmp838 & tmp840) | (tmp839 & tmp840);
  wire tmp842;
  assign tmp842 = 1'b0;
  wire tmp843;
  assign tmp843 = 1'b0;
  wire tmp844;
  assign tmp844 = 1'b0;
  wire tmp845;
  assign tmp845 = (tmp842 & tmp843) | (tmp842 & tmp844) | (tmp843 & tmp844);
  wire tmp846;
  assign tmp846 = (tmp837 & tmp841) | (tmp837 & tmp845) | (tmp841 & tmp845);
  wire tmp847;
  assign tmp847 = (tmp820 & tmp833) | (tmp820 & tmp846) | (tmp833 & tmp846);
  wire tmp848;
  assign tmp848 = (tmp767 & tmp807) | (tmp767 & tmp847) | (tmp807 & tmp847);
  wire tmp849;
  assign tmp849 = pi1;
  wire tmp850;
  assign tmp850 = 1'b1;
  wire tmp851;
  assign tmp851 = 1'b1;
  wire tmp852;
  assign tmp852 = (tmp849 & tmp850) | (tmp849 & tmp851) | (tmp850 & tmp851);
  wire tmp853;
  assign tmp853 = 1'b1;
  wire tmp854;
  assign tmp854 = 1'b0;
  wire tmp855;
  assign tmp855 = 1'b0;
  wire tmp856;
  assign tmp856 = (tmp853 & tmp854) | (tmp853 & tmp855) | (tmp854 & tmp855);
  wire tmp857;
  assign tmp857 = 1'b1;
  wire tmp858;
  assign tmp858 = 1'b0;
  wire tmp859;
  assign tmp859 = 1'b0;
  wire tmp860;
  assign tmp860 = (tmp857 & tmp858) | (tmp857 & tmp859) | (tmp858 & tmp859);
  wire tmp861;
  assign tmp861 = (tmp852 & tmp856) | (tmp852 & tmp860) | (tmp856 & tmp860);
  wire tmp862;
  assign tmp862 = 1'b1;
  wire tmp863;
  assign tmp863 = 1'b0;
  wire tmp864;
  assign tmp864 = 1'b0;
  wire tmp865;
  assign tmp865 = (tmp862 & tmp863) | (tmp862 & tmp864) | (tmp863 & tmp864);
  wire tmp866;
  assign tmp866 = 1'b0;
  wire tmp867;
  assign tmp867 = pi3;
  wire tmp868;
  assign tmp868 = 1'b0;
  wire tmp869;
  assign tmp869 = (tmp866 & tmp867) | (tmp866 & tmp868) | (tmp867 & tmp868);
  wire tmp870;
  assign tmp870 = 1'b0;
  wire tmp871;
  assign tmp871 = 1'b0;
  wire tmp872;
  assign tmp872 = 1'b0;
  wire tmp873;
  assign tmp873 = (tmp870 & tmp871) | (tmp870 & tmp872) | (tmp871 & tmp872);
  wire tmp874;
  assign tmp874 = (tmp865 & tmp869) | (tmp865 & tmp873) | (tmp869 & tmp873);
  wire tmp875;
  assign tmp875 = 1'b1;
  wire tmp876;
  assign tmp876 = 1'b0;
  wire tmp877;
  assign tmp877 = 1'b0;
  wire tmp878;
  assign tmp878 = (tmp875 & tmp876) | (tmp875 & tmp877) | (tmp876 & tmp877);
  wire tmp879;
  assign tmp879 = 1'b0;
  wire tmp880;
  assign tmp880 = 1'b0;
  wire tmp881;
  assign tmp881 = 1'b0;
  wire tmp882;
  assign tmp882 = (tmp879 & tmp880) | (tmp879 & tmp881) | (tmp880 & tmp881);
  wire tmp883;
  assign tmp883 = 1'b0;
  wire tmp884;
  assign tmp884 = 1'b0;
  wire tmp885;
  assign tmp885 = 1'b0;
  wire tmp886;
  assign tmp886 = (tmp883 & tmp884) | (tmp883 & tmp885) | (tmp884 & tmp885);
  wire tmp887;
  assign tmp887 = (tmp878 & tmp882) | (tmp878 & tmp886) | (tmp882 & tmp886);
  wire tmp888;
  assign tmp888 = (tmp861 & tmp874) | (tmp861 & tmp887) | (tmp874 & tmp887);
  wire tmp889;
  assign tmp889 = 1'b1;
  wire tmp890;
  assign tmp890 = 1'b0;
  wire tmp891;
  assign tmp891 = 1'b0;
  wire tmp892;
  assign tmp892 = (tmp889 & tmp890) | (tmp889 & tmp891) | (tmp890 & tmp891);
  wire tmp893;
  assign tmp893 = 1'b0;
  wire tmp894;
  assign tmp894 = pi3;
  wire tmp895;
  assign tmp895 = 1'b0;
  wire tmp896;
  assign tmp896 = (tmp893 & tmp894) | (tmp893 & tmp895) | (tmp894 & tmp895);
  wire tmp897;
  assign tmp897 = 1'b0;
  wire tmp898;
  assign tmp898 = 1'b0;
  wire tmp899;
  assign tmp899 = 1'b0;
  wire tmp900;
  assign tmp900 = (tmp897 & tmp898) | (tmp897 & tmp899) | (tmp898 & tmp899);
  wire tmp901;
  assign tmp901 = (tmp892 & tmp896) | (tmp892 & tmp900) | (tmp896 & tmp900);
  wire tmp902;
  assign tmp902 = 1'b0;
  wire tmp903;
  assign tmp903 = pi3;
  wire tmp904;
  assign tmp904 = 1'b0;
  wire tmp905;
  assign tmp905 = (tmp902 & tmp903) | (tmp902 & tmp904) | (tmp903 & tmp904);
  wire tmp906;
  assign tmp906 = pi3;
  wire tmp907;
  assign tmp907 = 1'b1;
  wire tmp908;
  assign tmp908 = 1'b0;
  wire tmp909;
  assign tmp909 = (tmp906 & tmp907) | (tmp906 & tmp908) | (tmp907 & tmp908);
  wire tmp910;
  assign tmp910 = 1'b0;
  wire tmp911;
  assign tmp911 = 1'b0;
  wire tmp912;
  assign tmp912 = 1'b0;
  wire tmp913;
  assign tmp913 = (tmp910 & tmp911) | (tmp910 & tmp912) | (tmp911 & tmp912);
  wire tmp914;
  assign tmp914 = (tmp905 & tmp909) | (tmp905 & tmp913) | (tmp909 & tmp913);
  wire tmp915;
  assign tmp915 = 1'b0;
  wire tmp916;
  assign tmp916 = 1'b0;
  wire tmp917;
  assign tmp917 = 1'b0;
  wire tmp918;
  assign tmp918 = (tmp915 & tmp916) | (tmp915 & tmp917) | (tmp916 & tmp917);
  wire tmp919;
  assign tmp919 = 1'b0;
  wire tmp920;
  assign tmp920 = 1'b0;
  wire tmp921;
  assign tmp921 = 1'b0;
  wire tmp922;
  assign tmp922 = (tmp919 & tmp920) | (tmp919 & tmp921) | (tmp920 & tmp921);
  wire tmp923;
  assign tmp923 = 1'b0;
  wire tmp924;
  assign tmp924 = 1'b0;
  wire tmp925;
  assign tmp925 = 1'b0;
  wire tmp926;
  assign tmp926 = (tmp923 & tmp924) | (tmp923 & tmp925) | (tmp924 & tmp925);
  wire tmp927;
  assign tmp927 = (tmp918 & tmp922) | (tmp918 & tmp926) | (tmp922 & tmp926);
  wire tmp928;
  assign tmp928 = (tmp901 & tmp914) | (tmp901 & tmp927) | (tmp914 & tmp927);
  wire tmp929;
  assign tmp929 = 1'b1;
  wire tmp930;
  assign tmp930 = 1'b0;
  wire tmp931;
  assign tmp931 = 1'b0;
  wire tmp932;
  assign tmp932 = (tmp929 & tmp930) | (tmp929 & tmp931) | (tmp930 & tmp931);
  wire tmp933;
  assign tmp933 = 1'b0;
  wire tmp934;
  assign tmp934 = 1'b0;
  wire tmp935;
  assign tmp935 = 1'b0;
  wire tmp936;
  assign tmp936 = (tmp933 & tmp934) | (tmp933 & tmp935) | (tmp934 & tmp935);
  wire tmp937;
  assign tmp937 = 1'b0;
  wire tmp938;
  assign tmp938 = 1'b0;
  wire tmp939;
  assign tmp939 = 1'b0;
  wire tmp940;
  assign tmp940 = (tmp937 & tmp938) | (tmp937 & tmp939) | (tmp938 & tmp939);
  wire tmp941;
  assign tmp941 = (tmp932 & tmp936) | (tmp932 & tmp940) | (tmp936 & tmp940);
  wire tmp942;
  assign tmp942 = 1'b0;
  wire tmp943;
  assign tmp943 = 1'b0;
  wire tmp944;
  assign tmp944 = 1'b0;
  wire tmp945;
  assign tmp945 = (tmp942 & tmp943) | (tmp942 & tmp944) | (tmp943 & tmp944);
  wire tmp946;
  assign tmp946 = 1'b0;
  wire tmp947;
  assign tmp947 = 1'b0;
  wire tmp948;
  assign tmp948 = 1'b0;
  wire tmp949;
  assign tmp949 = (tmp946 & tmp947) | (tmp946 & tmp948) | (tmp947 & tmp948);
  wire tmp950;
  assign tmp950 = 1'b0;
  wire tmp951;
  assign tmp951 = 1'b0;
  wire tmp952;
  assign tmp952 = 1'b0;
  wire tmp953;
  assign tmp953 = (tmp950 & tmp951) | (tmp950 & tmp952) | (tmp951 & tmp952);
  wire tmp954;
  assign tmp954 = (tmp945 & tmp949) | (tmp945 & tmp953) | (tmp949 & tmp953);
  wire tmp955;
  assign tmp955 = 1'b0;
  wire tmp956;
  assign tmp956 = 1'b0;
  wire tmp957;
  assign tmp957 = 1'b0;
  wire tmp958;
  assign tmp958 = (tmp955 & tmp956) | (tmp955 & tmp957) | (tmp956 & tmp957);
  wire tmp959;
  assign tmp959 = 1'b0;
  wire tmp960;
  assign tmp960 = 1'b0;
  wire tmp961;
  assign tmp961 = 1'b0;
  wire tmp962;
  assign tmp962 = (tmp959 & tmp960) | (tmp959 & tmp961) | (tmp960 & tmp961);
  wire tmp963;
  assign tmp963 = 1'b0;
  wire tmp964;
  assign tmp964 = 1'b0;
  wire tmp965;
  assign tmp965 = 1'b0;
  wire tmp966;
  assign tmp966 = (tmp963 & tmp964) | (tmp963 & tmp965) | (tmp964 & tmp965);
  wire tmp967;
  assign tmp967 = (tmp958 & tmp962) | (tmp958 & tmp966) | (tmp962 & tmp966);
  wire tmp968;
  assign tmp968 = (tmp941 & tmp954) | (tmp941 & tmp967) | (tmp954 & tmp967);
  wire tmp969;
  assign tmp969 = (tmp888 & tmp928) | (tmp888 & tmp968) | (tmp928 & tmp968);
  wire tmp970;
  assign tmp970 = pi4;
  wire tmp971;
  assign tmp971 = 1'b1;
  wire tmp972;
  assign tmp972 = 1'b0;
  wire tmp973;
  assign tmp973 = (tmp970 & tmp971) | (tmp970 & tmp972) | (tmp971 & tmp972);
  wire tmp974;
  assign tmp974 = 1'b1;
  wire tmp975;
  assign tmp975 = 1'b0;
  wire tmp976;
  assign tmp976 = 1'b0;
  wire tmp977;
  assign tmp977 = (tmp974 & tmp975) | (tmp974 & tmp976) | (tmp975 & tmp976);
  wire tmp978;
  assign tmp978 = 1'b0;
  wire tmp979;
  assign tmp979 = 1'b0;
  wire tmp980;
  assign tmp980 = 1'b0;
  wire tmp981;
  assign tmp981 = (tmp978 & tmp979) | (tmp978 & tmp980) | (tmp979 & tmp980);
  wire tmp982;
  assign tmp982 = (tmp973 & tmp977) | (tmp973 & tmp981) | (tmp977 & tmp981);
  wire tmp983;
  assign tmp983 = 1'b1;
  wire tmp984;
  assign tmp984 = 1'b0;
  wire tmp985;
  assign tmp985 = 1'b0;
  wire tmp986;
  assign tmp986 = (tmp983 & tmp984) | (tmp983 & tmp985) | (tmp984 & tmp985);
  wire tmp987;
  assign tmp987 = 1'b0;
  wire tmp988;
  assign tmp988 = 1'b0;
  wire tmp989;
  assign tmp989 = 1'b0;
  wire tmp990;
  assign tmp990 = (tmp987 & tmp988) | (tmp987 & tmp989) | (tmp988 & tmp989);
  wire tmp991;
  assign tmp991 = 1'b0;
  wire tmp992;
  assign tmp992 = 1'b0;
  wire tmp993;
  assign tmp993 = 1'b0;
  wire tmp994;
  assign tmp994 = (tmp991 & tmp992) | (tmp991 & tmp993) | (tmp992 & tmp993);
  wire tmp995;
  assign tmp995 = (tmp986 & tmp990) | (tmp986 & tmp994) | (tmp990 & tmp994);
  wire tmp996;
  assign tmp996 = 1'b0;
  wire tmp997;
  assign tmp997 = 1'b0;
  wire tmp998;
  assign tmp998 = 1'b0;
  wire tmp999;
  assign tmp999 = (tmp996 & tmp997) | (tmp996 & tmp998) | (tmp997 & tmp998);
  wire tmp1000;
  assign tmp1000 = 1'b0;
  wire tmp1001;
  assign tmp1001 = 1'b0;
  wire tmp1002;
  assign tmp1002 = 1'b0;
  wire tmp1003;
  assign tmp1003 = (tmp1000 & tmp1001) | (tmp1000 & tmp1002) | (tmp1001 & tmp1002);
  wire tmp1004;
  assign tmp1004 = 1'b0;
  wire tmp1005;
  assign tmp1005 = 1'b0;
  wire tmp1006;
  assign tmp1006 = 1'b0;
  wire tmp1007;
  assign tmp1007 = (tmp1004 & tmp1005) | (tmp1004 & tmp1006) | (tmp1005 & tmp1006);
  wire tmp1008;
  assign tmp1008 = (tmp999 & tmp1003) | (tmp999 & tmp1007) | (tmp1003 & tmp1007);
  wire tmp1009;
  assign tmp1009 = (tmp982 & tmp995) | (tmp982 & tmp1008) | (tmp995 & tmp1008);
  wire tmp1010;
  assign tmp1010 = 1'b1;
  wire tmp1011;
  assign tmp1011 = 1'b0;
  wire tmp1012;
  assign tmp1012 = 1'b0;
  wire tmp1013;
  assign tmp1013 = (tmp1010 & tmp1011) | (tmp1010 & tmp1012) | (tmp1011 & tmp1012);
  wire tmp1014;
  assign tmp1014 = 1'b0;
  wire tmp1015;
  assign tmp1015 = 1'b0;
  wire tmp1016;
  assign tmp1016 = 1'b0;
  wire tmp1017;
  assign tmp1017 = (tmp1014 & tmp1015) | (tmp1014 & tmp1016) | (tmp1015 & tmp1016);
  wire tmp1018;
  assign tmp1018 = 1'b0;
  wire tmp1019;
  assign tmp1019 = 1'b0;
  wire tmp1020;
  assign tmp1020 = 1'b0;
  wire tmp1021;
  assign tmp1021 = (tmp1018 & tmp1019) | (tmp1018 & tmp1020) | (tmp1019 & tmp1020);
  wire tmp1022;
  assign tmp1022 = (tmp1013 & tmp1017) | (tmp1013 & tmp1021) | (tmp1017 & tmp1021);
  wire tmp1023;
  assign tmp1023 = 1'b0;
  wire tmp1024;
  assign tmp1024 = 1'b0;
  wire tmp1025;
  assign tmp1025 = 1'b0;
  wire tmp1026;
  assign tmp1026 = (tmp1023 & tmp1024) | (tmp1023 & tmp1025) | (tmp1024 & tmp1025);
  wire tmp1027;
  assign tmp1027 = 1'b0;
  wire tmp1028;
  assign tmp1028 = 1'b0;
  wire tmp1029;
  assign tmp1029 = 1'b0;
  wire tmp1030;
  assign tmp1030 = (tmp1027 & tmp1028) | (tmp1027 & tmp1029) | (tmp1028 & tmp1029);
  wire tmp1031;
  assign tmp1031 = 1'b0;
  wire tmp1032;
  assign tmp1032 = 1'b0;
  wire tmp1033;
  assign tmp1033 = 1'b0;
  wire tmp1034;
  assign tmp1034 = (tmp1031 & tmp1032) | (tmp1031 & tmp1033) | (tmp1032 & tmp1033);
  wire tmp1035;
  assign tmp1035 = (tmp1026 & tmp1030) | (tmp1026 & tmp1034) | (tmp1030 & tmp1034);
  wire tmp1036;
  assign tmp1036 = 1'b0;
  wire tmp1037;
  assign tmp1037 = 1'b0;
  wire tmp1038;
  assign tmp1038 = 1'b0;
  wire tmp1039;
  assign tmp1039 = (tmp1036 & tmp1037) | (tmp1036 & tmp1038) | (tmp1037 & tmp1038);
  wire tmp1040;
  assign tmp1040 = 1'b0;
  wire tmp1041;
  assign tmp1041 = 1'b0;
  wire tmp1042;
  assign tmp1042 = 1'b0;
  wire tmp1043;
  assign tmp1043 = (tmp1040 & tmp1041) | (tmp1040 & tmp1042) | (tmp1041 & tmp1042);
  wire tmp1044;
  assign tmp1044 = 1'b0;
  wire tmp1045;
  assign tmp1045 = 1'b0;
  wire tmp1046;
  assign tmp1046 = 1'b0;
  wire tmp1047;
  assign tmp1047 = (tmp1044 & tmp1045) | (tmp1044 & tmp1046) | (tmp1045 & tmp1046);
  wire tmp1048;
  assign tmp1048 = (tmp1039 & tmp1043) | (tmp1039 & tmp1047) | (tmp1043 & tmp1047);
  wire tmp1049;
  assign tmp1049 = (tmp1022 & tmp1035) | (tmp1022 & tmp1048) | (tmp1035 & tmp1048);
  wire tmp1050;
  assign tmp1050 = 1'b0;
  wire tmp1051;
  assign tmp1051 = 1'b0;
  wire tmp1052;
  assign tmp1052 = 1'b0;
  wire tmp1053;
  assign tmp1053 = (tmp1050 & tmp1051) | (tmp1050 & tmp1052) | (tmp1051 & tmp1052);
  wire tmp1054;
  assign tmp1054 = 1'b0;
  wire tmp1055;
  assign tmp1055 = 1'b0;
  wire tmp1056;
  assign tmp1056 = 1'b0;
  wire tmp1057;
  assign tmp1057 = (tmp1054 & tmp1055) | (tmp1054 & tmp1056) | (tmp1055 & tmp1056);
  wire tmp1058;
  assign tmp1058 = 1'b0;
  wire tmp1059;
  assign tmp1059 = 1'b0;
  wire tmp1060;
  assign tmp1060 = 1'b0;
  wire tmp1061;
  assign tmp1061 = (tmp1058 & tmp1059) | (tmp1058 & tmp1060) | (tmp1059 & tmp1060);
  wire tmp1062;
  assign tmp1062 = (tmp1053 & tmp1057) | (tmp1053 & tmp1061) | (tmp1057 & tmp1061);
  wire tmp1063;
  assign tmp1063 = 1'b0;
  wire tmp1064;
  assign tmp1064 = 1'b0;
  wire tmp1065;
  assign tmp1065 = 1'b0;
  wire tmp1066;
  assign tmp1066 = (tmp1063 & tmp1064) | (tmp1063 & tmp1065) | (tmp1064 & tmp1065);
  wire tmp1067;
  assign tmp1067 = 1'b0;
  wire tmp1068;
  assign tmp1068 = 1'b0;
  wire tmp1069;
  assign tmp1069 = 1'b0;
  wire tmp1070;
  assign tmp1070 = (tmp1067 & tmp1068) | (tmp1067 & tmp1069) | (tmp1068 & tmp1069);
  wire tmp1071;
  assign tmp1071 = 1'b0;
  wire tmp1072;
  assign tmp1072 = 1'b0;
  wire tmp1073;
  assign tmp1073 = 1'b0;
  wire tmp1074;
  assign tmp1074 = (tmp1071 & tmp1072) | (tmp1071 & tmp1073) | (tmp1072 & tmp1073);
  wire tmp1075;
  assign tmp1075 = (tmp1066 & tmp1070) | (tmp1066 & tmp1074) | (tmp1070 & tmp1074);
  wire tmp1076;
  assign tmp1076 = 1'b0;
  wire tmp1077;
  assign tmp1077 = 1'b0;
  wire tmp1078;
  assign tmp1078 = 1'b0;
  wire tmp1079;
  assign tmp1079 = (tmp1076 & tmp1077) | (tmp1076 & tmp1078) | (tmp1077 & tmp1078);
  wire tmp1080;
  assign tmp1080 = 1'b0;
  wire tmp1081;
  assign tmp1081 = 1'b0;
  wire tmp1082;
  assign tmp1082 = 1'b0;
  wire tmp1083;
  assign tmp1083 = (tmp1080 & tmp1081) | (tmp1080 & tmp1082) | (tmp1081 & tmp1082);
  wire tmp1084;
  assign tmp1084 = 1'b0;
  wire tmp1085;
  assign tmp1085 = 1'b0;
  wire tmp1086;
  assign tmp1086 = 1'b0;
  wire tmp1087;
  assign tmp1087 = (tmp1084 & tmp1085) | (tmp1084 & tmp1086) | (tmp1085 & tmp1086);
  wire tmp1088;
  assign tmp1088 = (tmp1079 & tmp1083) | (tmp1079 & tmp1087) | (tmp1083 & tmp1087);
  wire tmp1089;
  assign tmp1089 = (tmp1062 & tmp1075) | (tmp1062 & tmp1088) | (tmp1075 & tmp1088);
  wire tmp1090;
  assign tmp1090 = (tmp1009 & tmp1049) | (tmp1009 & tmp1089) | (tmp1049 & tmp1089);
  wire tmp1091;
  assign tmp1091 = (tmp848 & tmp969) | (tmp848 & tmp1090) | (tmp969 & tmp1090);
  wire tmp1092;
  assign tmp1092 = (tmp363 & tmp727) | (tmp363 & tmp1091) | (tmp727 & tmp1091);
  assign po0 = tmp1092;
endmodule // test_4
