module test_inv( pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, po0 );
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
  output po0;
  wire tmp0;
  assign tmp0 = pi0;
  wire tmp1;
  assign tmp1 = pi1;
  wire tmp2;
  assign tmp2 = 1'b0;
  wire tmp3;
  assign tmp3 = (tmp0 & tmp1) | (tmp0 & tmp2) | (tmp1 & tmp2);
  wire tmp4;
  assign tmp4 = pi1;
  wire tmp5;
  assign tmp5 = pi2;
  wire tmp6;
  assign tmp6 = 1'b0;
  wire tmp7;
  assign tmp7 = (tmp4 & tmp5) | (tmp4 & tmp6) | (tmp5 & tmp6);
  wire tmp8;
  assign tmp8 = 1'b0;
  wire tmp9;
  assign tmp9 = 1'b0;
  wire tmp10;
  assign tmp10 = 1'b0;
  wire tmp11;
  assign tmp11 = (tmp8 & tmp9) | (tmp8 & tmp10) | (tmp9 & tmp10);
  wire tmp12;
  assign tmp12 = (tmp3 & tmp7) | (tmp3 & tmp11) | (tmp7 & tmp11);
  wire tmp13;
  assign tmp13 = pi1;
  wire tmp14;
  assign tmp14 = pi2;
  wire tmp15;
  assign tmp15 = 1'b0;
  wire tmp16;
  assign tmp16 = (tmp13 & tmp14) | (tmp13 & tmp15) | (tmp14 & tmp15);
  wire tmp17;
  assign tmp17 = pi2;
  wire tmp18;
  assign tmp18 = pi3;
  wire tmp19;
  assign tmp19 = 1'b0;
  wire tmp20;
  assign tmp20 = (tmp17 & tmp18) | (tmp17 & tmp19) | (tmp18 & tmp19);
  wire tmp21;
  assign tmp21 = 1'b0;
  wire tmp22;
  assign tmp22 = 1'b0;
  wire tmp23;
  assign tmp23 = 1'b0;
  wire tmp24;
  assign tmp24 = (tmp21 & tmp22) | (tmp21 & tmp23) | (tmp22 & tmp23);
  wire tmp25;
  assign tmp25 = (tmp16 & tmp20) | (tmp16 & tmp24) | (tmp20 & tmp24);
  wire tmp26;
  assign tmp26 = 1'b0;
  wire tmp27;
  assign tmp27 = 1'b0;
  wire tmp28;
  assign tmp28 = 1'b0;
  wire tmp29;
  assign tmp29 = (tmp26 & tmp27) | (tmp26 & tmp28) | (tmp27 & tmp28);
  wire tmp30;
  assign tmp30 = 1'b0;
  wire tmp31;
  assign tmp31 = 1'b0;
  wire tmp32;
  assign tmp32 = 1'b0;
  wire tmp33;
  assign tmp33 = (tmp30 & tmp31) | (tmp30 & tmp32) | (tmp31 & tmp32);
  wire tmp34;
  assign tmp34 = 1'b0;
  wire tmp35;
  assign tmp35 = 1'b0;
  wire tmp36;
  assign tmp36 = 1'b0;
  wire tmp37;
  assign tmp37 = (tmp34 & tmp35) | (tmp34 & tmp36) | (tmp35 & tmp36);
  wire tmp38;
  assign tmp38 = (tmp29 & tmp33) | (tmp29 & tmp37) | (tmp33 & tmp37);
  wire tmp39;
  assign tmp39 = (tmp12 & tmp25) | (tmp12 & tmp38) | (tmp25 & tmp38);
  wire tmp40;
  assign tmp40 = pi1;
  wire tmp41;
  assign tmp41 = pi2;
  wire tmp42;
  assign tmp42 = 1'b0;
  wire tmp43;
  assign tmp43 = (tmp40 & tmp41) | (tmp40 & tmp42) | (tmp41 & tmp42);
  wire tmp44;
  assign tmp44 = pi2;
  wire tmp45;
  assign tmp45 = pi3;
  wire tmp46;
  assign tmp46 = 1'b0;
  wire tmp47;
  assign tmp47 = (tmp44 & tmp45) | (tmp44 & tmp46) | (tmp45 & tmp46);
  wire tmp48;
  assign tmp48 = 1'b0;
  wire tmp49;
  assign tmp49 = 1'b0;
  wire tmp50;
  assign tmp50 = 1'b0;
  wire tmp51;
  assign tmp51 = (tmp48 & tmp49) | (tmp48 & tmp50) | (tmp49 & tmp50);
  wire tmp52;
  assign tmp52 = (tmp43 & tmp47) | (tmp43 & tmp51) | (tmp47 & tmp51);
  wire tmp53;
  assign tmp53 = pi2;
  wire tmp54;
  assign tmp54 = pi3;
  wire tmp55;
  assign tmp55 = 1'b0;
  wire tmp56;
  assign tmp56 = (tmp53 & tmp54) | (tmp53 & tmp55) | (tmp54 & tmp55);
  wire tmp57;
  assign tmp57 = pi3;
  wire tmp58;
  assign tmp58 = 1'b1;
  wire tmp59;
  assign tmp59 = 1'b0;
  wire tmp60;
  assign tmp60 = (tmp57 & tmp58) | (tmp57 & tmp59) | (tmp58 & tmp59);
  wire tmp61;
  assign tmp61 = 1'b0;
  wire tmp62;
  assign tmp62 = 1'b0;
  wire tmp63;
  assign tmp63 = 1'b0;
  wire tmp64;
  assign tmp64 = (tmp61 & tmp62) | (tmp61 & tmp63) | (tmp62 & tmp63);
  wire tmp65;
  assign tmp65 = (tmp56 & tmp60) | (tmp56 & tmp64) | (tmp60 & tmp64);
  wire tmp66;
  assign tmp66 = 1'b0;
  wire tmp67;
  assign tmp67 = 1'b0;
  wire tmp68;
  assign tmp68 = 1'b0;
  wire tmp69;
  assign tmp69 = (tmp66 & tmp67) | (tmp66 & tmp68) | (tmp67 & tmp68);
  wire tmp70;
  assign tmp70 = 1'b0;
  wire tmp71;
  assign tmp71 = 1'b0;
  wire tmp72;
  assign tmp72 = 1'b0;
  wire tmp73;
  assign tmp73 = (tmp70 & tmp71) | (tmp70 & tmp72) | (tmp71 & tmp72);
  wire tmp74;
  assign tmp74 = 1'b0;
  wire tmp75;
  assign tmp75 = 1'b0;
  wire tmp76;
  assign tmp76 = 1'b0;
  wire tmp77;
  assign tmp77 = (tmp74 & tmp75) | (tmp74 & tmp76) | (tmp75 & tmp76);
  wire tmp78;
  assign tmp78 = (tmp69 & tmp73) | (tmp69 & tmp77) | (tmp73 & tmp77);
  wire tmp79;
  assign tmp79 = (tmp52 & tmp65) | (tmp52 & tmp78) | (tmp65 & tmp78);
  wire tmp80;
  assign tmp80 = 1'b0;
  wire tmp81;
  assign tmp81 = 1'b0;
  wire tmp82;
  assign tmp82 = 1'b0;
  wire tmp83;
  assign tmp83 = (tmp80 & tmp81) | (tmp80 & tmp82) | (tmp81 & tmp82);
  wire tmp84;
  assign tmp84 = 1'b0;
  wire tmp85;
  assign tmp85 = 1'b0;
  wire tmp86;
  assign tmp86 = 1'b0;
  wire tmp87;
  assign tmp87 = (tmp84 & tmp85) | (tmp84 & tmp86) | (tmp85 & tmp86);
  wire tmp88;
  assign tmp88 = 1'b0;
  wire tmp89;
  assign tmp89 = 1'b0;
  wire tmp90;
  assign tmp90 = 1'b0;
  wire tmp91;
  assign tmp91 = (tmp88 & tmp89) | (tmp88 & tmp90) | (tmp89 & tmp90);
  wire tmp92;
  assign tmp92 = (tmp83 & tmp87) | (tmp83 & tmp91) | (tmp87 & tmp91);
  wire tmp93;
  assign tmp93 = 1'b0;
  wire tmp94;
  assign tmp94 = 1'b0;
  wire tmp95;
  assign tmp95 = 1'b0;
  wire tmp96;
  assign tmp96 = (tmp93 & tmp94) | (tmp93 & tmp95) | (tmp94 & tmp95);
  wire tmp97;
  assign tmp97 = 1'b0;
  wire tmp98;
  assign tmp98 = 1'b0;
  wire tmp99;
  assign tmp99 = 1'b0;
  wire tmp100;
  assign tmp100 = (tmp97 & tmp98) | (tmp97 & tmp99) | (tmp98 & tmp99);
  wire tmp101;
  assign tmp101 = 1'b0;
  wire tmp102;
  assign tmp102 = 1'b0;
  wire tmp103;
  assign tmp103 = 1'b0;
  wire tmp104;
  assign tmp104 = (tmp101 & tmp102) | (tmp101 & tmp103) | (tmp102 & tmp103);
  wire tmp105;
  assign tmp105 = (tmp96 & tmp100) | (tmp96 & tmp104) | (tmp100 & tmp104);
  wire tmp106;
  assign tmp106 = 1'b0;
  wire tmp107;
  assign tmp107 = 1'b0;
  wire tmp108;
  assign tmp108 = 1'b0;
  wire tmp109;
  assign tmp109 = (tmp106 & tmp107) | (tmp106 & tmp108) | (tmp107 & tmp108);
  wire tmp110;
  assign tmp110 = 1'b0;
  wire tmp111;
  assign tmp111 = 1'b0;
  wire tmp112;
  assign tmp112 = 1'b0;
  wire tmp113;
  assign tmp113 = (tmp110 & tmp111) | (tmp110 & tmp112) | (tmp111 & tmp112);
  wire tmp114;
  assign tmp114 = 1'b0;
  wire tmp115;
  assign tmp115 = 1'b0;
  wire tmp116;
  assign tmp116 = 1'b0;
  wire tmp117;
  assign tmp117 = (tmp114 & tmp115) | (tmp114 & tmp116) | (tmp115 & tmp116);
  wire tmp118;
  assign tmp118 = (tmp109 & tmp113) | (tmp109 & tmp117) | (tmp113 & tmp117);
  wire tmp119;
  assign tmp119 = (tmp92 & tmp105) | (tmp92 & tmp118) | (tmp105 & tmp118);
  wire tmp120;
  assign tmp120 = (tmp39 & tmp79) | (tmp39 & tmp119) | (tmp79 & tmp119);
  wire tmp121;
  assign tmp121 = pi1;
  wire tmp122;
  assign tmp122 = pi2;
  wire tmp123;
  assign tmp123 = 1'b0;
  wire tmp124;
  assign tmp124 = (tmp121 & tmp122) | (tmp121 & tmp123) | (tmp122 & tmp123);
  wire tmp125;
  assign tmp125 = pi2;
  wire tmp126;
  assign tmp126 = pi3;
  wire tmp127;
  assign tmp127 = 1'b0;
  wire tmp128;
  assign tmp128 = (tmp125 & tmp126) | (tmp125 & tmp127) | (tmp126 & tmp127);
  wire tmp129;
  assign tmp129 = 1'b0;
  wire tmp130;
  assign tmp130 = 1'b0;
  wire tmp131;
  assign tmp131 = 1'b0;
  wire tmp132;
  assign tmp132 = (tmp129 & tmp130) | (tmp129 & tmp131) | (tmp130 & tmp131);
  wire tmp133;
  assign tmp133 = (tmp124 & tmp128) | (tmp124 & tmp132) | (tmp128 & tmp132);
  wire tmp134;
  assign tmp134 = pi2;
  wire tmp135;
  assign tmp135 = pi3;
  wire tmp136;
  assign tmp136 = 1'b0;
  wire tmp137;
  assign tmp137 = (tmp134 & tmp135) | (tmp134 & tmp136) | (tmp135 & tmp136);
  wire tmp138;
  assign tmp138 = pi3;
  wire tmp139;
  assign tmp139 = 1'b1;
  wire tmp140;
  assign tmp140 = 1'b0;
  wire tmp141;
  assign tmp141 = (tmp138 & tmp139) | (tmp138 & tmp140) | (tmp139 & tmp140);
  wire tmp142;
  assign tmp142 = 1'b0;
  wire tmp143;
  assign tmp143 = 1'b0;
  wire tmp144;
  assign tmp144 = 1'b0;
  wire tmp145;
  assign tmp145 = (tmp142 & tmp143) | (tmp142 & tmp144) | (tmp143 & tmp144);
  wire tmp146;
  assign tmp146 = (tmp137 & tmp141) | (tmp137 & tmp145) | (tmp141 & tmp145);
  wire tmp147;
  assign tmp147 = 1'b0;
  wire tmp148;
  assign tmp148 = 1'b0;
  wire tmp149;
  assign tmp149 = 1'b0;
  wire tmp150;
  assign tmp150 = (tmp147 & tmp148) | (tmp147 & tmp149) | (tmp148 & tmp149);
  wire tmp151;
  assign tmp151 = 1'b0;
  wire tmp152;
  assign tmp152 = 1'b0;
  wire tmp153;
  assign tmp153 = 1'b0;
  wire tmp154;
  assign tmp154 = (tmp151 & tmp152) | (tmp151 & tmp153) | (tmp152 & tmp153);
  wire tmp155;
  assign tmp155 = 1'b0;
  wire tmp156;
  assign tmp156 = 1'b0;
  wire tmp157;
  assign tmp157 = 1'b0;
  wire tmp158;
  assign tmp158 = (tmp155 & tmp156) | (tmp155 & tmp157) | (tmp156 & tmp157);
  wire tmp159;
  assign tmp159 = (tmp150 & tmp154) | (tmp150 & tmp158) | (tmp154 & tmp158);
  wire tmp160;
  assign tmp160 = (tmp133 & tmp146) | (tmp133 & tmp159) | (tmp146 & tmp159);
  wire tmp161;
  assign tmp161 = pi2;
  wire tmp162;
  assign tmp162 = pi3;
  wire tmp163;
  assign tmp163 = 1'b0;
  wire tmp164;
  assign tmp164 = (tmp161 & tmp162) | (tmp161 & tmp163) | (tmp162 & tmp163);
  wire tmp165;
  assign tmp165 = pi3;
  wire tmp166;
  assign tmp166 = 1'b1;
  wire tmp167;
  assign tmp167 = 1'b0;
  wire tmp168;
  assign tmp168 = (tmp165 & tmp166) | (tmp165 & tmp167) | (tmp166 & tmp167);
  wire tmp169;
  assign tmp169 = 1'b0;
  wire tmp170;
  assign tmp170 = 1'b0;
  wire tmp171;
  assign tmp171 = 1'b0;
  wire tmp172;
  assign tmp172 = (tmp169 & tmp170) | (tmp169 & tmp171) | (tmp170 & tmp171);
  wire tmp173;
  assign tmp173 = (tmp164 & tmp168) | (tmp164 & tmp172) | (tmp168 & tmp172);
  wire tmp174;
  assign tmp174 = pi3;
  wire tmp175;
  assign tmp175 = 1'b1;
  wire tmp176;
  assign tmp176 = 1'b0;
  wire tmp177;
  assign tmp177 = (tmp174 & tmp175) | (tmp174 & tmp176) | (tmp175 & tmp176);
  wire tmp178;
  assign tmp178 = 1'b1;
  wire tmp179;
  assign tmp179 = 1'b1;
  wire tmp180;
  assign tmp180 = 1'b1;
  wire tmp181;
  assign tmp181 = (tmp178 & tmp179) | (tmp178 & tmp180) | (tmp179 & tmp180);
  wire tmp182;
  assign tmp182 = 1'b0;
  wire tmp183;
  assign tmp183 = 1'b1;
  wire tmp184;
  assign tmp184 = 1'b0;
  wire tmp185;
  assign tmp185 = (tmp182 & tmp183) | (tmp182 & tmp184) | (tmp183 & tmp184);
  wire tmp186;
  assign tmp186 = (tmp177 & tmp181) | (tmp177 & tmp185) | (tmp181 & tmp185);
  wire tmp187;
  assign tmp187 = 1'b0;
  wire tmp188;
  assign tmp188 = 1'b0;
  wire tmp189;
  assign tmp189 = 1'b0;
  wire tmp190;
  assign tmp190 = (tmp187 & tmp188) | (tmp187 & tmp189) | (tmp188 & tmp189);
  wire tmp191;
  assign tmp191 = 1'b0;
  wire tmp192;
  assign tmp192 = 1'b1;
  wire tmp193;
  assign tmp193 = 1'b0;
  wire tmp194;
  assign tmp194 = (tmp191 & tmp192) | (tmp191 & tmp193) | (tmp192 & tmp193);
  wire tmp195;
  assign tmp195 = 1'b0;
  wire tmp196;
  assign tmp196 = 1'b0;
  wire tmp197;
  assign tmp197 = 1'b0;
  wire tmp198;
  assign tmp198 = (tmp195 & tmp196) | (tmp195 & tmp197) | (tmp196 & tmp197);
  wire tmp199;
  assign tmp199 = (tmp190 & tmp194) | (tmp190 & tmp198) | (tmp194 & tmp198);
  wire tmp200;
  assign tmp200 = (tmp173 & tmp186) | (tmp173 & tmp199) | (tmp186 & tmp199);
  wire tmp201;
  assign tmp201 = 1'b0;
  wire tmp202;
  assign tmp202 = 1'b0;
  wire tmp203;
  assign tmp203 = 1'b0;
  wire tmp204;
  assign tmp204 = (tmp201 & tmp202) | (tmp201 & tmp203) | (tmp202 & tmp203);
  wire tmp205;
  assign tmp205 = 1'b0;
  wire tmp206;
  assign tmp206 = 1'b0;
  wire tmp207;
  assign tmp207 = 1'b0;
  wire tmp208;
  assign tmp208 = (tmp205 & tmp206) | (tmp205 & tmp207) | (tmp206 & tmp207);
  wire tmp209;
  assign tmp209 = 1'b0;
  wire tmp210;
  assign tmp210 = 1'b0;
  wire tmp211;
  assign tmp211 = 1'b0;
  wire tmp212;
  assign tmp212 = (tmp209 & tmp210) | (tmp209 & tmp211) | (tmp210 & tmp211);
  wire tmp213;
  assign tmp213 = (tmp204 & tmp208) | (tmp204 & tmp212) | (tmp208 & tmp212);
  wire tmp214;
  assign tmp214 = 1'b0;
  wire tmp215;
  assign tmp215 = 1'b0;
  wire tmp216;
  assign tmp216 = 1'b0;
  wire tmp217;
  assign tmp217 = (tmp214 & tmp215) | (tmp214 & tmp216) | (tmp215 & tmp216);
  wire tmp218;
  assign tmp218 = 1'b0;
  wire tmp219;
  assign tmp219 = 1'b1;
  wire tmp220;
  assign tmp220 = 1'b0;
  wire tmp221;
  assign tmp221 = (tmp218 & tmp219) | (tmp218 & tmp220) | (tmp219 & tmp220);
  wire tmp222;
  assign tmp222 = 1'b0;
  wire tmp223;
  assign tmp223 = 1'b0;
  wire tmp224;
  assign tmp224 = 1'b0;
  wire tmp225;
  assign tmp225 = (tmp222 & tmp223) | (tmp222 & tmp224) | (tmp223 & tmp224);
  wire tmp226;
  assign tmp226 = (tmp217 & tmp221) | (tmp217 & tmp225) | (tmp221 & tmp225);
  wire tmp227;
  assign tmp227 = 1'b0;
  wire tmp228;
  assign tmp228 = 1'b0;
  wire tmp229;
  assign tmp229 = 1'b0;
  wire tmp230;
  assign tmp230 = (tmp227 & tmp228) | (tmp227 & tmp229) | (tmp228 & tmp229);
  wire tmp231;
  assign tmp231 = 1'b0;
  wire tmp232;
  assign tmp232 = 1'b0;
  wire tmp233;
  assign tmp233 = 1'b0;
  wire tmp234;
  assign tmp234 = (tmp231 & tmp232) | (tmp231 & tmp233) | (tmp232 & tmp233);
  wire tmp235;
  assign tmp235 = 1'b0;
  wire tmp236;
  assign tmp236 = 1'b0;
  wire tmp237;
  assign tmp237 = 1'b0;
  wire tmp238;
  assign tmp238 = (tmp235 & tmp236) | (tmp235 & tmp237) | (tmp236 & tmp237);
  wire tmp239;
  assign tmp239 = (tmp230 & tmp234) | (tmp230 & tmp238) | (tmp234 & tmp238);
  wire tmp240;
  assign tmp240 = (tmp213 & tmp226) | (tmp213 & tmp239) | (tmp226 & tmp239);
  wire tmp241;
  assign tmp241 = (tmp160 & tmp200) | (tmp160 & tmp240) | (tmp200 & tmp240);
  wire tmp242;
  assign tmp242 = 1'b0;
  wire tmp243;
  assign tmp243 = 1'b0;
  wire tmp244;
  assign tmp244 = 1'b0;
  wire tmp245;
  assign tmp245 = (tmp242 & tmp243) | (tmp242 & tmp244) | (tmp243 & tmp244);
  wire tmp246;
  assign tmp246 = 1'b0;
  wire tmp247;
  assign tmp247 = 1'b0;
  wire tmp248;
  assign tmp248 = 1'b0;
  wire tmp249;
  assign tmp249 = (tmp246 & tmp247) | (tmp246 & tmp248) | (tmp247 & tmp248);
  wire tmp250;
  assign tmp250 = 1'b0;
  wire tmp251;
  assign tmp251 = 1'b0;
  wire tmp252;
  assign tmp252 = 1'b0;
  wire tmp253;
  assign tmp253 = (tmp250 & tmp251) | (tmp250 & tmp252) | (tmp251 & tmp252);
  wire tmp254;
  assign tmp254 = (tmp245 & tmp249) | (tmp245 & tmp253) | (tmp249 & tmp253);
  wire tmp255;
  assign tmp255 = 1'b0;
  wire tmp256;
  assign tmp256 = 1'b0;
  wire tmp257;
  assign tmp257 = 1'b0;
  wire tmp258;
  assign tmp258 = (tmp255 & tmp256) | (tmp255 & tmp257) | (tmp256 & tmp257);
  wire tmp259;
  assign tmp259 = 1'b0;
  wire tmp260;
  assign tmp260 = 1'b0;
  wire tmp261;
  assign tmp261 = 1'b0;
  wire tmp262;
  assign tmp262 = (tmp259 & tmp260) | (tmp259 & tmp261) | (tmp260 & tmp261);
  wire tmp263;
  assign tmp263 = 1'b0;
  wire tmp264;
  assign tmp264 = 1'b0;
  wire tmp265;
  assign tmp265 = 1'b0;
  wire tmp266;
  assign tmp266 = (tmp263 & tmp264) | (tmp263 & tmp265) | (tmp264 & tmp265);
  wire tmp267;
  assign tmp267 = (tmp258 & tmp262) | (tmp258 & tmp266) | (tmp262 & tmp266);
  wire tmp268;
  assign tmp268 = 1'b0;
  wire tmp269;
  assign tmp269 = 1'b0;
  wire tmp270;
  assign tmp270 = 1'b0;
  wire tmp271;
  assign tmp271 = (tmp268 & tmp269) | (tmp268 & tmp270) | (tmp269 & tmp270);
  wire tmp272;
  assign tmp272 = 1'b0;
  wire tmp273;
  assign tmp273 = 1'b0;
  wire tmp274;
  assign tmp274 = 1'b0;
  wire tmp275;
  assign tmp275 = (tmp272 & tmp273) | (tmp272 & tmp274) | (tmp273 & tmp274);
  wire tmp276;
  assign tmp276 = 1'b0;
  wire tmp277;
  assign tmp277 = 1'b0;
  wire tmp278;
  assign tmp278 = 1'b0;
  wire tmp279;
  assign tmp279 = (tmp276 & tmp277) | (tmp276 & tmp278) | (tmp277 & tmp278);
  wire tmp280;
  assign tmp280 = (tmp271 & tmp275) | (tmp271 & tmp279) | (tmp275 & tmp279);
  wire tmp281;
  assign tmp281 = (tmp254 & tmp267) | (tmp254 & tmp280) | (tmp267 & tmp280);
  wire tmp282;
  assign tmp282 = 1'b0;
  wire tmp283;
  assign tmp283 = 1'b0;
  wire tmp284;
  assign tmp284 = 1'b0;
  wire tmp285;
  assign tmp285 = (tmp282 & tmp283) | (tmp282 & tmp284) | (tmp283 & tmp284);
  wire tmp286;
  assign tmp286 = 1'b0;
  wire tmp287;
  assign tmp287 = 1'b0;
  wire tmp288;
  assign tmp288 = 1'b0;
  wire tmp289;
  assign tmp289 = (tmp286 & tmp287) | (tmp286 & tmp288) | (tmp287 & tmp288);
  wire tmp290;
  assign tmp290 = 1'b0;
  wire tmp291;
  assign tmp291 = 1'b0;
  wire tmp292;
  assign tmp292 = 1'b0;
  wire tmp293;
  assign tmp293 = (tmp290 & tmp291) | (tmp290 & tmp292) | (tmp291 & tmp292);
  wire tmp294;
  assign tmp294 = (tmp285 & tmp289) | (tmp285 & tmp293) | (tmp289 & tmp293);
  wire tmp295;
  assign tmp295 = 1'b0;
  wire tmp296;
  assign tmp296 = 1'b0;
  wire tmp297;
  assign tmp297 = 1'b0;
  wire tmp298;
  assign tmp298 = (tmp295 & tmp296) | (tmp295 & tmp297) | (tmp296 & tmp297);
  wire tmp299;
  assign tmp299 = 1'b0;
  wire tmp300;
  assign tmp300 = 1'b1;
  wire tmp301;
  assign tmp301 = 1'b0;
  wire tmp302;
  assign tmp302 = (tmp299 & tmp300) | (tmp299 & tmp301) | (tmp300 & tmp301);
  wire tmp303;
  assign tmp303 = 1'b0;
  wire tmp304;
  assign tmp304 = 1'b0;
  wire tmp305;
  assign tmp305 = 1'b0;
  wire tmp306;
  assign tmp306 = (tmp303 & tmp304) | (tmp303 & tmp305) | (tmp304 & tmp305);
  wire tmp307;
  assign tmp307 = (tmp298 & tmp302) | (tmp298 & tmp306) | (tmp302 & tmp306);
  wire tmp308;
  assign tmp308 = 1'b0;
  wire tmp309;
  assign tmp309 = 1'b0;
  wire tmp310;
  assign tmp310 = 1'b0;
  wire tmp311;
  assign tmp311 = (tmp308 & tmp309) | (tmp308 & tmp310) | (tmp309 & tmp310);
  wire tmp312;
  assign tmp312 = 1'b0;
  wire tmp313;
  assign tmp313 = 1'b0;
  wire tmp314;
  assign tmp314 = 1'b0;
  wire tmp315;
  assign tmp315 = (tmp312 & tmp313) | (tmp312 & tmp314) | (tmp313 & tmp314);
  wire tmp316;
  assign tmp316 = 1'b0;
  wire tmp317;
  assign tmp317 = 1'b0;
  wire tmp318;
  assign tmp318 = 1'b0;
  wire tmp319;
  assign tmp319 = (tmp316 & tmp317) | (tmp316 & tmp318) | (tmp317 & tmp318);
  wire tmp320;
  assign tmp320 = (tmp311 & tmp315) | (tmp311 & tmp319) | (tmp315 & tmp319);
  wire tmp321;
  assign tmp321 = (tmp294 & tmp307) | (tmp294 & tmp320) | (tmp307 & tmp320);
  wire tmp322;
  assign tmp322 = 1'b0;
  wire tmp323;
  assign tmp323 = 1'b0;
  wire tmp324;
  assign tmp324 = 1'b0;
  wire tmp325;
  assign tmp325 = (tmp322 & tmp323) | (tmp322 & tmp324) | (tmp323 & tmp324);
  wire tmp326;
  assign tmp326 = 1'b0;
  wire tmp327;
  assign tmp327 = 1'b0;
  wire tmp328;
  assign tmp328 = 1'b0;
  wire tmp329;
  assign tmp329 = (tmp326 & tmp327) | (tmp326 & tmp328) | (tmp327 & tmp328);
  wire tmp330;
  assign tmp330 = 1'b0;
  wire tmp331;
  assign tmp331 = 1'b0;
  wire tmp332;
  assign tmp332 = 1'b0;
  wire tmp333;
  assign tmp333 = (tmp330 & tmp331) | (tmp330 & tmp332) | (tmp331 & tmp332);
  wire tmp334;
  assign tmp334 = (tmp325 & tmp329) | (tmp325 & tmp333) | (tmp329 & tmp333);
  wire tmp335;
  assign tmp335 = 1'b0;
  wire tmp336;
  assign tmp336 = 1'b0;
  wire tmp337;
  assign tmp337 = 1'b0;
  wire tmp338;
  assign tmp338 = (tmp335 & tmp336) | (tmp335 & tmp337) | (tmp336 & tmp337);
  wire tmp339;
  assign tmp339 = 1'b0;
  wire tmp340;
  assign tmp340 = 1'b0;
  wire tmp341;
  assign tmp341 = 1'b0;
  wire tmp342;
  assign tmp342 = (tmp339 & tmp340) | (tmp339 & tmp341) | (tmp340 & tmp341);
  wire tmp343;
  assign tmp343 = 1'b0;
  wire tmp344;
  assign tmp344 = 1'b0;
  wire tmp345;
  assign tmp345 = 1'b0;
  wire tmp346;
  assign tmp346 = (tmp343 & tmp344) | (tmp343 & tmp345) | (tmp344 & tmp345);
  wire tmp347;
  assign tmp347 = (tmp338 & tmp342) | (tmp338 & tmp346) | (tmp342 & tmp346);
  wire tmp348;
  assign tmp348 = 1'b0;
  wire tmp349;
  assign tmp349 = 1'b0;
  wire tmp350;
  assign tmp350 = 1'b0;
  wire tmp351;
  assign tmp351 = (tmp348 & tmp349) | (tmp348 & tmp350) | (tmp349 & tmp350);
  wire tmp352;
  assign tmp352 = 1'b0;
  wire tmp353;
  assign tmp353 = 1'b0;
  wire tmp354;
  assign tmp354 = 1'b0;
  wire tmp355;
  assign tmp355 = (tmp352 & tmp353) | (tmp352 & tmp354) | (tmp353 & tmp354);
  wire tmp356;
  assign tmp356 = 1'b0;
  wire tmp357;
  assign tmp357 = 1'b0;
  wire tmp358;
  assign tmp358 = 1'b0;
  wire tmp359;
  assign tmp359 = (tmp356 & tmp357) | (tmp356 & tmp358) | (tmp357 & tmp358);
  wire tmp360;
  assign tmp360 = (tmp351 & tmp355) | (tmp351 & tmp359) | (tmp355 & tmp359);
  wire tmp361;
  assign tmp361 = (tmp334 & tmp347) | (tmp334 & tmp360) | (tmp347 & tmp360);
  wire tmp362;
  assign tmp362 = (tmp281 & tmp321) | (tmp281 & tmp361) | (tmp321 & tmp361);
  wire tmp363;
  assign tmp363 = (tmp120 & tmp241) | (tmp120 & tmp362) | (tmp241 & tmp362);
  wire tmp364;
  assign tmp364 = pi1;
  wire tmp365;
  assign tmp365 = pi2;
  wire tmp366;
  assign tmp366 = 1'b0;
  wire tmp367;
  assign tmp367 = (tmp364 & tmp365) | (tmp364 & tmp366) | (tmp365 & tmp366);
  wire tmp368;
  assign tmp368 = pi2;
  wire tmp369;
  assign tmp369 = pi3;
  wire tmp370;
  assign tmp370 = 1'b0;
  wire tmp371;
  assign tmp371 = (tmp368 & tmp369) | (tmp368 & tmp370) | (tmp369 & tmp370);
  wire tmp372;
  assign tmp372 = 1'b0;
  wire tmp373;
  assign tmp373 = 1'b0;
  wire tmp374;
  assign tmp374 = 1'b0;
  wire tmp375;
  assign tmp375 = (tmp372 & tmp373) | (tmp372 & tmp374) | (tmp373 & tmp374);
  wire tmp376;
  assign tmp376 = (tmp367 & tmp371) | (tmp367 & tmp375) | (tmp371 & tmp375);
  wire tmp377;
  assign tmp377 = pi2;
  wire tmp378;
  assign tmp378 = pi3;
  wire tmp379;
  assign tmp379 = 1'b0;
  wire tmp380;
  assign tmp380 = (tmp377 & tmp378) | (tmp377 & tmp379) | (tmp378 & tmp379);
  wire tmp381;
  assign tmp381 = pi3;
  wire tmp382;
  assign tmp382 = 1'b1;
  wire tmp383;
  assign tmp383 = 1'b0;
  wire tmp384;
  assign tmp384 = (tmp381 & tmp382) | (tmp381 & tmp383) | (tmp382 & tmp383);
  wire tmp385;
  assign tmp385 = 1'b0;
  wire tmp386;
  assign tmp386 = 1'b0;
  wire tmp387;
  assign tmp387 = 1'b0;
  wire tmp388;
  assign tmp388 = (tmp385 & tmp386) | (tmp385 & tmp387) | (tmp386 & tmp387);
  wire tmp389;
  assign tmp389 = (tmp380 & tmp384) | (tmp380 & tmp388) | (tmp384 & tmp388);
  wire tmp390;
  assign tmp390 = 1'b0;
  wire tmp391;
  assign tmp391 = 1'b0;
  wire tmp392;
  assign tmp392 = 1'b0;
  wire tmp393;
  assign tmp393 = (tmp390 & tmp391) | (tmp390 & tmp392) | (tmp391 & tmp392);
  wire tmp394;
  assign tmp394 = 1'b0;
  wire tmp395;
  assign tmp395 = 1'b0;
  wire tmp396;
  assign tmp396 = 1'b0;
  wire tmp397;
  assign tmp397 = (tmp394 & tmp395) | (tmp394 & tmp396) | (tmp395 & tmp396);
  wire tmp398;
  assign tmp398 = 1'b0;
  wire tmp399;
  assign tmp399 = 1'b0;
  wire tmp400;
  assign tmp400 = 1'b0;
  wire tmp401;
  assign tmp401 = (tmp398 & tmp399) | (tmp398 & tmp400) | (tmp399 & tmp400);
  wire tmp402;
  assign tmp402 = (tmp393 & tmp397) | (tmp393 & tmp401) | (tmp397 & tmp401);
  wire tmp403;
  assign tmp403 = (tmp376 & tmp389) | (tmp376 & tmp402) | (tmp389 & tmp402);
  wire tmp404;
  assign tmp404 = pi2;
  wire tmp405;
  assign tmp405 = pi3;
  wire tmp406;
  assign tmp406 = 1'b0;
  wire tmp407;
  assign tmp407 = (tmp404 & tmp405) | (tmp404 & tmp406) | (tmp405 & tmp406);
  wire tmp408;
  assign tmp408 = pi3;
  wire tmp409;
  assign tmp409 = 1'b1;
  wire tmp410;
  assign tmp410 = 1'b0;
  wire tmp411;
  assign tmp411 = (tmp408 & tmp409) | (tmp408 & tmp410) | (tmp409 & tmp410);
  wire tmp412;
  assign tmp412 = 1'b0;
  wire tmp413;
  assign tmp413 = 1'b0;
  wire tmp414;
  assign tmp414 = 1'b0;
  wire tmp415;
  assign tmp415 = (tmp412 & tmp413) | (tmp412 & tmp414) | (tmp413 & tmp414);
  wire tmp416;
  assign tmp416 = (tmp407 & tmp411) | (tmp407 & tmp415) | (tmp411 & tmp415);
  wire tmp417;
  assign tmp417 = pi3;
  wire tmp418;
  assign tmp418 = 1'b1;
  wire tmp419;
  assign tmp419 = 1'b0;
  wire tmp420;
  assign tmp420 = (tmp417 & tmp418) | (tmp417 & tmp419) | (tmp418 & tmp419);
  wire tmp421;
  assign tmp421 = 1'b1;
  wire tmp422;
  assign tmp422 = 1'b1;
  wire tmp423;
  assign tmp423 = 1'b1;
  wire tmp424;
  assign tmp424 = (tmp421 & tmp422) | (tmp421 & tmp423) | (tmp422 & tmp423);
  wire tmp425;
  assign tmp425 = 1'b0;
  wire tmp426;
  assign tmp426 = 1'b1;
  wire tmp427;
  assign tmp427 = 1'b0;
  wire tmp428;
  assign tmp428 = (tmp425 & tmp426) | (tmp425 & tmp427) | (tmp426 & tmp427);
  wire tmp429;
  assign tmp429 = (tmp420 & tmp424) | (tmp420 & tmp428) | (tmp424 & tmp428);
  wire tmp430;
  assign tmp430 = 1'b0;
  wire tmp431;
  assign tmp431 = 1'b0;
  wire tmp432;
  assign tmp432 = 1'b0;
  wire tmp433;
  assign tmp433 = (tmp430 & tmp431) | (tmp430 & tmp432) | (tmp431 & tmp432);
  wire tmp434;
  assign tmp434 = 1'b0;
  wire tmp435;
  assign tmp435 = 1'b1;
  wire tmp436;
  assign tmp436 = 1'b0;
  wire tmp437;
  assign tmp437 = (tmp434 & tmp435) | (tmp434 & tmp436) | (tmp435 & tmp436);
  wire tmp438;
  assign tmp438 = 1'b0;
  wire tmp439;
  assign tmp439 = 1'b0;
  wire tmp440;
  assign tmp440 = 1'b0;
  wire tmp441;
  assign tmp441 = (tmp438 & tmp439) | (tmp438 & tmp440) | (tmp439 & tmp440);
  wire tmp442;
  assign tmp442 = (tmp433 & tmp437) | (tmp433 & tmp441) | (tmp437 & tmp441);
  wire tmp443;
  assign tmp443 = (tmp416 & tmp429) | (tmp416 & tmp442) | (tmp429 & tmp442);
  wire tmp444;
  assign tmp444 = 1'b0;
  wire tmp445;
  assign tmp445 = 1'b0;
  wire tmp446;
  assign tmp446 = 1'b0;
  wire tmp447;
  assign tmp447 = (tmp444 & tmp445) | (tmp444 & tmp446) | (tmp445 & tmp446);
  wire tmp448;
  assign tmp448 = 1'b0;
  wire tmp449;
  assign tmp449 = 1'b0;
  wire tmp450;
  assign tmp450 = 1'b0;
  wire tmp451;
  assign tmp451 = (tmp448 & tmp449) | (tmp448 & tmp450) | (tmp449 & tmp450);
  wire tmp452;
  assign tmp452 = 1'b0;
  wire tmp453;
  assign tmp453 = 1'b0;
  wire tmp454;
  assign tmp454 = 1'b0;
  wire tmp455;
  assign tmp455 = (tmp452 & tmp453) | (tmp452 & tmp454) | (tmp453 & tmp454);
  wire tmp456;
  assign tmp456 = (tmp447 & tmp451) | (tmp447 & tmp455) | (tmp451 & tmp455);
  wire tmp457;
  assign tmp457 = 1'b0;
  wire tmp458;
  assign tmp458 = 1'b0;
  wire tmp459;
  assign tmp459 = 1'b0;
  wire tmp460;
  assign tmp460 = (tmp457 & tmp458) | (tmp457 & tmp459) | (tmp458 & tmp459);
  wire tmp461;
  assign tmp461 = 1'b0;
  wire tmp462;
  assign tmp462 = 1'b1;
  wire tmp463;
  assign tmp463 = 1'b0;
  wire tmp464;
  assign tmp464 = (tmp461 & tmp462) | (tmp461 & tmp463) | (tmp462 & tmp463);
  wire tmp465;
  assign tmp465 = 1'b0;
  wire tmp466;
  assign tmp466 = 1'b0;
  wire tmp467;
  assign tmp467 = 1'b0;
  wire tmp468;
  assign tmp468 = (tmp465 & tmp466) | (tmp465 & tmp467) | (tmp466 & tmp467);
  wire tmp469;
  assign tmp469 = (tmp460 & tmp464) | (tmp460 & tmp468) | (tmp464 & tmp468);
  wire tmp470;
  assign tmp470 = 1'b0;
  wire tmp471;
  assign tmp471 = 1'b0;
  wire tmp472;
  assign tmp472 = 1'b0;
  wire tmp473;
  assign tmp473 = (tmp470 & tmp471) | (tmp470 & tmp472) | (tmp471 & tmp472);
  wire tmp474;
  assign tmp474 = 1'b0;
  wire tmp475;
  assign tmp475 = 1'b0;
  wire tmp476;
  assign tmp476 = 1'b0;
  wire tmp477;
  assign tmp477 = (tmp474 & tmp475) | (tmp474 & tmp476) | (tmp475 & tmp476);
  wire tmp478;
  assign tmp478 = 1'b0;
  wire tmp479;
  assign tmp479 = 1'b0;
  wire tmp480;
  assign tmp480 = 1'b0;
  wire tmp481;
  assign tmp481 = (tmp478 & tmp479) | (tmp478 & tmp480) | (tmp479 & tmp480);
  wire tmp482;
  assign tmp482 = (tmp473 & tmp477) | (tmp473 & tmp481) | (tmp477 & tmp481);
  wire tmp483;
  assign tmp483 = (tmp456 & tmp469) | (tmp456 & tmp482) | (tmp469 & tmp482);
  wire tmp484;
  assign tmp484 = (tmp403 & tmp443) | (tmp403 & tmp483) | (tmp443 & tmp483);
  wire tmp485;
  assign tmp485 = pi2;
  wire tmp486;
  assign tmp486 = pi3;
  wire tmp487;
  assign tmp487 = 1'b0;
  wire tmp488;
  assign tmp488 = (tmp485 & tmp486) | (tmp485 & tmp487) | (tmp486 & tmp487);
  wire tmp489;
  assign tmp489 = pi3;
  wire tmp490;
  assign tmp490 = 1'b1;
  wire tmp491;
  assign tmp491 = 1'b0;
  wire tmp492;
  assign tmp492 = (tmp489 & tmp490) | (tmp489 & tmp491) | (tmp490 & tmp491);
  wire tmp493;
  assign tmp493 = 1'b0;
  wire tmp494;
  assign tmp494 = 1'b0;
  wire tmp495;
  assign tmp495 = 1'b0;
  wire tmp496;
  assign tmp496 = (tmp493 & tmp494) | (tmp493 & tmp495) | (tmp494 & tmp495);
  wire tmp497;
  assign tmp497 = (tmp488 & tmp492) | (tmp488 & tmp496) | (tmp492 & tmp496);
  wire tmp498;
  assign tmp498 = pi3;
  wire tmp499;
  assign tmp499 = 1'b1;
  wire tmp500;
  assign tmp500 = 1'b0;
  wire tmp501;
  assign tmp501 = (tmp498 & tmp499) | (tmp498 & tmp500) | (tmp499 & tmp500);
  wire tmp502;
  assign tmp502 = 1'b1;
  wire tmp503;
  assign tmp503 = 1'b1;
  wire tmp504;
  assign tmp504 = 1'b1;
  wire tmp505;
  assign tmp505 = (tmp502 & tmp503) | (tmp502 & tmp504) | (tmp503 & tmp504);
  wire tmp506;
  assign tmp506 = 1'b0;
  wire tmp507;
  assign tmp507 = 1'b1;
  wire tmp508;
  assign tmp508 = 1'b0;
  wire tmp509;
  assign tmp509 = (tmp506 & tmp507) | (tmp506 & tmp508) | (tmp507 & tmp508);
  wire tmp510;
  assign tmp510 = (tmp501 & tmp505) | (tmp501 & tmp509) | (tmp505 & tmp509);
  wire tmp511;
  assign tmp511 = 1'b0;
  wire tmp512;
  assign tmp512 = 1'b0;
  wire tmp513;
  assign tmp513 = 1'b0;
  wire tmp514;
  assign tmp514 = (tmp511 & tmp512) | (tmp511 & tmp513) | (tmp512 & tmp513);
  wire tmp515;
  assign tmp515 = 1'b0;
  wire tmp516;
  assign tmp516 = 1'b1;
  wire tmp517;
  assign tmp517 = 1'b0;
  wire tmp518;
  assign tmp518 = (tmp515 & tmp516) | (tmp515 & tmp517) | (tmp516 & tmp517);
  wire tmp519;
  assign tmp519 = 1'b0;
  wire tmp520;
  assign tmp520 = 1'b0;
  wire tmp521;
  assign tmp521 = 1'b0;
  wire tmp522;
  assign tmp522 = (tmp519 & tmp520) | (tmp519 & tmp521) | (tmp520 & tmp521);
  wire tmp523;
  assign tmp523 = (tmp514 & tmp518) | (tmp514 & tmp522) | (tmp518 & tmp522);
  wire tmp524;
  assign tmp524 = (tmp497 & tmp510) | (tmp497 & tmp523) | (tmp510 & tmp523);
  wire tmp525;
  assign tmp525 = pi3;
  wire tmp526;
  assign tmp526 = 1'b1;
  wire tmp527;
  assign tmp527 = 1'b0;
  wire tmp528;
  assign tmp528 = (tmp525 & tmp526) | (tmp525 & tmp527) | (tmp526 & tmp527);
  wire tmp529;
  assign tmp529 = 1'b1;
  wire tmp530;
  assign tmp530 = 1'b1;
  wire tmp531;
  assign tmp531 = 1'b1;
  wire tmp532;
  assign tmp532 = (tmp529 & tmp530) | (tmp529 & tmp531) | (tmp530 & tmp531);
  wire tmp533;
  assign tmp533 = 1'b0;
  wire tmp534;
  assign tmp534 = 1'b1;
  wire tmp535;
  assign tmp535 = 1'b0;
  wire tmp536;
  assign tmp536 = (tmp533 & tmp534) | (tmp533 & tmp535) | (tmp534 & tmp535);
  wire tmp537;
  assign tmp537 = (tmp528 & tmp532) | (tmp528 & tmp536) | (tmp532 & tmp536);
  wire tmp538;
  assign tmp538 = 1'b1;
  wire tmp539;
  assign tmp539 = 1'b1;
  wire tmp540;
  assign tmp540 = 1'b1;
  wire tmp541;
  assign tmp541 = (tmp538 & tmp539) | (tmp538 & tmp540) | (tmp539 & tmp540);
  wire tmp542;
  assign tmp542 = 1'b1;
  wire tmp543;
  assign tmp543 = 1'b1;
  wire tmp544;
  assign tmp544 = 1'b1;
  wire tmp545;
  assign tmp545 = (tmp542 & tmp543) | (tmp542 & tmp544) | (tmp543 & tmp544);
  wire tmp546;
  assign tmp546 = 1'b1;
  wire tmp547;
  assign tmp547 = 1'b1;
  wire tmp548;
  assign tmp548 = 1'b1;
  wire tmp549;
  assign tmp549 = (tmp546 & tmp547) | (tmp546 & tmp548) | (tmp547 & tmp548);
  wire tmp550;
  assign tmp550 = (tmp541 & tmp545) | (tmp541 & tmp549) | (tmp545 & tmp549);
  wire tmp551;
  assign tmp551 = 1'b0;
  wire tmp552;
  assign tmp552 = 1'b1;
  wire tmp553;
  assign tmp553 = 1'b0;
  wire tmp554;
  assign tmp554 = (tmp551 & tmp552) | (tmp551 & tmp553) | (tmp552 & tmp553);
  wire tmp555;
  assign tmp555 = 1'b1;
  wire tmp556;
  assign tmp556 = 1'b1;
  wire tmp557;
  assign tmp557 = 1'b1;
  wire tmp558;
  assign tmp558 = (tmp555 & tmp556) | (tmp555 & tmp557) | (tmp556 & tmp557);
  wire tmp559;
  assign tmp559 = 1'b0;
  wire tmp560;
  assign tmp560 = 1'b1;
  wire tmp561;
  assign tmp561 = 1'b0;
  wire tmp562;
  assign tmp562 = (tmp559 & tmp560) | (tmp559 & tmp561) | (tmp560 & tmp561);
  wire tmp563;
  assign tmp563 = (tmp554 & tmp558) | (tmp554 & tmp562) | (tmp558 & tmp562);
  wire tmp564;
  assign tmp564 = (tmp537 & tmp550) | (tmp537 & tmp563) | (tmp550 & tmp563);
  wire tmp565;
  assign tmp565 = 1'b0;
  wire tmp566;
  assign tmp566 = 1'b0;
  wire tmp567;
  assign tmp567 = 1'b0;
  wire tmp568;
  assign tmp568 = (tmp565 & tmp566) | (tmp565 & tmp567) | (tmp566 & tmp567);
  wire tmp569;
  assign tmp569 = 1'b0;
  wire tmp570;
  assign tmp570 = 1'b1;
  wire tmp571;
  assign tmp571 = 1'b0;
  wire tmp572;
  assign tmp572 = (tmp569 & tmp570) | (tmp569 & tmp571) | (tmp570 & tmp571);
  wire tmp573;
  assign tmp573 = 1'b0;
  wire tmp574;
  assign tmp574 = 1'b0;
  wire tmp575;
  assign tmp575 = 1'b0;
  wire tmp576;
  assign tmp576 = (tmp573 & tmp574) | (tmp573 & tmp575) | (tmp574 & tmp575);
  wire tmp577;
  assign tmp577 = (tmp568 & tmp572) | (tmp568 & tmp576) | (tmp572 & tmp576);
  wire tmp578;
  assign tmp578 = 1'b0;
  wire tmp579;
  assign tmp579 = 1'b1;
  wire tmp580;
  assign tmp580 = 1'b0;
  wire tmp581;
  assign tmp581 = (tmp578 & tmp579) | (tmp578 & tmp580) | (tmp579 & tmp580);
  wire tmp582;
  assign tmp582 = 1'b1;
  wire tmp583;
  assign tmp583 = 1'b1;
  wire tmp584;
  assign tmp584 = 1'b1;
  wire tmp585;
  assign tmp585 = (tmp582 & tmp583) | (tmp582 & tmp584) | (tmp583 & tmp584);
  wire tmp586;
  assign tmp586 = 1'b0;
  wire tmp587;
  assign tmp587 = 1'b1;
  wire tmp588;
  assign tmp588 = 1'b0;
  wire tmp589;
  assign tmp589 = (tmp586 & tmp587) | (tmp586 & tmp588) | (tmp587 & tmp588);
  wire tmp590;
  assign tmp590 = (tmp581 & tmp585) | (tmp581 & tmp589) | (tmp585 & tmp589);
  wire tmp591;
  assign tmp591 = 1'b0;
  wire tmp592;
  assign tmp592 = 1'b0;
  wire tmp593;
  assign tmp593 = 1'b0;
  wire tmp594;
  assign tmp594 = (tmp591 & tmp592) | (tmp591 & tmp593) | (tmp592 & tmp593);
  wire tmp595;
  assign tmp595 = 1'b0;
  wire tmp596;
  assign tmp596 = 1'b1;
  wire tmp597;
  assign tmp597 = 1'b0;
  wire tmp598;
  assign tmp598 = (tmp595 & tmp596) | (tmp595 & tmp597) | (tmp596 & tmp597);
  wire tmp599;
  assign tmp599 = 1'b0;
  wire tmp600;
  assign tmp600 = 1'b0;
  wire tmp601;
  assign tmp601 = 1'b0;
  wire tmp602;
  assign tmp602 = (tmp599 & tmp600) | (tmp599 & tmp601) | (tmp600 & tmp601);
  wire tmp603;
  assign tmp603 = (tmp594 & tmp598) | (tmp594 & tmp602) | (tmp598 & tmp602);
  wire tmp604;
  assign tmp604 = (tmp577 & tmp590) | (tmp577 & tmp603) | (tmp590 & tmp603);
  wire tmp605;
  assign tmp605 = (tmp524 & tmp564) | (tmp524 & tmp604) | (tmp564 & tmp604);
  wire tmp606;
  assign tmp606 = 1'b0;
  wire tmp607;
  assign tmp607 = 1'b0;
  wire tmp608;
  assign tmp608 = 1'b0;
  wire tmp609;
  assign tmp609 = (tmp606 & tmp607) | (tmp606 & tmp608) | (tmp607 & tmp608);
  wire tmp610;
  assign tmp610 = 1'b0;
  wire tmp611;
  assign tmp611 = 1'b0;
  wire tmp612;
  assign tmp612 = 1'b0;
  wire tmp613;
  assign tmp613 = (tmp610 & tmp611) | (tmp610 & tmp612) | (tmp611 & tmp612);
  wire tmp614;
  assign tmp614 = 1'b0;
  wire tmp615;
  assign tmp615 = 1'b0;
  wire tmp616;
  assign tmp616 = 1'b0;
  wire tmp617;
  assign tmp617 = (tmp614 & tmp615) | (tmp614 & tmp616) | (tmp615 & tmp616);
  wire tmp618;
  assign tmp618 = (tmp609 & tmp613) | (tmp609 & tmp617) | (tmp613 & tmp617);
  wire tmp619;
  assign tmp619 = 1'b0;
  wire tmp620;
  assign tmp620 = 1'b0;
  wire tmp621;
  assign tmp621 = 1'b0;
  wire tmp622;
  assign tmp622 = (tmp619 & tmp620) | (tmp619 & tmp621) | (tmp620 & tmp621);
  wire tmp623;
  assign tmp623 = 1'b0;
  wire tmp624;
  assign tmp624 = 1'b1;
  wire tmp625;
  assign tmp625 = 1'b0;
  wire tmp626;
  assign tmp626 = (tmp623 & tmp624) | (tmp623 & tmp625) | (tmp624 & tmp625);
  wire tmp627;
  assign tmp627 = 1'b0;
  wire tmp628;
  assign tmp628 = 1'b0;
  wire tmp629;
  assign tmp629 = 1'b0;
  wire tmp630;
  assign tmp630 = (tmp627 & tmp628) | (tmp627 & tmp629) | (tmp628 & tmp629);
  wire tmp631;
  assign tmp631 = (tmp622 & tmp626) | (tmp622 & tmp630) | (tmp626 & tmp630);
  wire tmp632;
  assign tmp632 = 1'b0;
  wire tmp633;
  assign tmp633 = 1'b0;
  wire tmp634;
  assign tmp634 = 1'b0;
  wire tmp635;
  assign tmp635 = (tmp632 & tmp633) | (tmp632 & tmp634) | (tmp633 & tmp634);
  wire tmp636;
  assign tmp636 = 1'b0;
  wire tmp637;
  assign tmp637 = 1'b0;
  wire tmp638;
  assign tmp638 = 1'b0;
  wire tmp639;
  assign tmp639 = (tmp636 & tmp637) | (tmp636 & tmp638) | (tmp637 & tmp638);
  wire tmp640;
  assign tmp640 = 1'b0;
  wire tmp641;
  assign tmp641 = 1'b0;
  wire tmp642;
  assign tmp642 = 1'b0;
  wire tmp643;
  assign tmp643 = (tmp640 & tmp641) | (tmp640 & tmp642) | (tmp641 & tmp642);
  wire tmp644;
  assign tmp644 = (tmp635 & tmp639) | (tmp635 & tmp643) | (tmp639 & tmp643);
  wire tmp645;
  assign tmp645 = (tmp618 & tmp631) | (tmp618 & tmp644) | (tmp631 & tmp644);
  wire tmp646;
  assign tmp646 = 1'b0;
  wire tmp647;
  assign tmp647 = 1'b0;
  wire tmp648;
  assign tmp648 = 1'b0;
  wire tmp649;
  assign tmp649 = (tmp646 & tmp647) | (tmp646 & tmp648) | (tmp647 & tmp648);
  wire tmp650;
  assign tmp650 = 1'b0;
  wire tmp651;
  assign tmp651 = 1'b1;
  wire tmp652;
  assign tmp652 = 1'b0;
  wire tmp653;
  assign tmp653 = (tmp650 & tmp651) | (tmp650 & tmp652) | (tmp651 & tmp652);
  wire tmp654;
  assign tmp654 = 1'b0;
  wire tmp655;
  assign tmp655 = 1'b0;
  wire tmp656;
  assign tmp656 = 1'b0;
  wire tmp657;
  assign tmp657 = (tmp654 & tmp655) | (tmp654 & tmp656) | (tmp655 & tmp656);
  wire tmp658;
  assign tmp658 = (tmp649 & tmp653) | (tmp649 & tmp657) | (tmp653 & tmp657);
  wire tmp659;
  assign tmp659 = 1'b0;
  wire tmp660;
  assign tmp660 = 1'b1;
  wire tmp661;
  assign tmp661 = 1'b0;
  wire tmp662;
  assign tmp662 = (tmp659 & tmp660) | (tmp659 & tmp661) | (tmp660 & tmp661);
  wire tmp663;
  assign tmp663 = 1'b1;
  wire tmp664;
  assign tmp664 = 1'b1;
  wire tmp665;
  assign tmp665 = 1'b1;
  wire tmp666;
  assign tmp666 = (tmp663 & tmp664) | (tmp663 & tmp665) | (tmp664 & tmp665);
  wire tmp667;
  assign tmp667 = 1'b0;
  wire tmp668;
  assign tmp668 = 1'b1;
  wire tmp669;
  assign tmp669 = 1'b0;
  wire tmp670;
  assign tmp670 = (tmp667 & tmp668) | (tmp667 & tmp669) | (tmp668 & tmp669);
  wire tmp671;
  assign tmp671 = (tmp662 & tmp666) | (tmp662 & tmp670) | (tmp666 & tmp670);
  wire tmp672;
  assign tmp672 = 1'b0;
  wire tmp673;
  assign tmp673 = 1'b0;
  wire tmp674;
  assign tmp674 = 1'b0;
  wire tmp675;
  assign tmp675 = (tmp672 & tmp673) | (tmp672 & tmp674) | (tmp673 & tmp674);
  wire tmp676;
  assign tmp676 = 1'b0;
  wire tmp677;
  assign tmp677 = 1'b1;
  wire tmp678;
  assign tmp678 = 1'b0;
  wire tmp679;
  assign tmp679 = (tmp676 & tmp677) | (tmp676 & tmp678) | (tmp677 & tmp678);
  wire tmp680;
  assign tmp680 = 1'b0;
  wire tmp681;
  assign tmp681 = 1'b0;
  wire tmp682;
  assign tmp682 = 1'b0;
  wire tmp683;
  assign tmp683 = (tmp680 & tmp681) | (tmp680 & tmp682) | (tmp681 & tmp682);
  wire tmp684;
  assign tmp684 = (tmp675 & tmp679) | (tmp675 & tmp683) | (tmp679 & tmp683);
  wire tmp685;
  assign tmp685 = (tmp658 & tmp671) | (tmp658 & tmp684) | (tmp671 & tmp684);
  wire tmp686;
  assign tmp686 = 1'b0;
  wire tmp687;
  assign tmp687 = 1'b0;
  wire tmp688;
  assign tmp688 = 1'b0;
  wire tmp689;
  assign tmp689 = (tmp686 & tmp687) | (tmp686 & tmp688) | (tmp687 & tmp688);
  wire tmp690;
  assign tmp690 = 1'b0;
  wire tmp691;
  assign tmp691 = 1'b0;
  wire tmp692;
  assign tmp692 = 1'b0;
  wire tmp693;
  assign tmp693 = (tmp690 & tmp691) | (tmp690 & tmp692) | (tmp691 & tmp692);
  wire tmp694;
  assign tmp694 = 1'b0;
  wire tmp695;
  assign tmp695 = 1'b0;
  wire tmp696;
  assign tmp696 = 1'b0;
  wire tmp697;
  assign tmp697 = (tmp694 & tmp695) | (tmp694 & tmp696) | (tmp695 & tmp696);
  wire tmp698;
  assign tmp698 = (tmp689 & tmp693) | (tmp689 & tmp697) | (tmp693 & tmp697);
  wire tmp699;
  assign tmp699 = 1'b0;
  wire tmp700;
  assign tmp700 = 1'b0;
  wire tmp701;
  assign tmp701 = 1'b0;
  wire tmp702;
  assign tmp702 = (tmp699 & tmp700) | (tmp699 & tmp701) | (tmp700 & tmp701);
  wire tmp703;
  assign tmp703 = 1'b0;
  wire tmp704;
  assign tmp704 = 1'b1;
  wire tmp705;
  assign tmp705 = 1'b0;
  wire tmp706;
  assign tmp706 = (tmp703 & tmp704) | (tmp703 & tmp705) | (tmp704 & tmp705);
  wire tmp707;
  assign tmp707 = 1'b0;
  wire tmp708;
  assign tmp708 = 1'b0;
  wire tmp709;
  assign tmp709 = 1'b0;
  wire tmp710;
  assign tmp710 = (tmp707 & tmp708) | (tmp707 & tmp709) | (tmp708 & tmp709);
  wire tmp711;
  assign tmp711 = (tmp702 & tmp706) | (tmp702 & tmp710) | (tmp706 & tmp710);
  wire tmp712;
  assign tmp712 = 1'b0;
  wire tmp713;
  assign tmp713 = 1'b0;
  wire tmp714;
  assign tmp714 = 1'b0;
  wire tmp715;
  assign tmp715 = (tmp712 & tmp713) | (tmp712 & tmp714) | (tmp713 & tmp714);
  wire tmp716;
  assign tmp716 = 1'b0;
  wire tmp717;
  assign tmp717 = 1'b0;
  wire tmp718;
  assign tmp718 = 1'b0;
  wire tmp719;
  assign tmp719 = (tmp716 & tmp717) | (tmp716 & tmp718) | (tmp717 & tmp718);
  wire tmp720;
  assign tmp720 = 1'b0;
  wire tmp721;
  assign tmp721 = 1'b0;
  wire tmp722;
  assign tmp722 = 1'b0;
  wire tmp723;
  assign tmp723 = (tmp720 & tmp721) | (tmp720 & tmp722) | (tmp721 & tmp722);
  wire tmp724;
  assign tmp724 = (tmp715 & tmp719) | (tmp715 & tmp723) | (tmp719 & tmp723);
  wire tmp725;
  assign tmp725 = (tmp698 & tmp711) | (tmp698 & tmp724) | (tmp711 & tmp724);
  wire tmp726;
  assign tmp726 = (tmp645 & tmp685) | (tmp645 & tmp725) | (tmp685 & tmp725);
  wire tmp727;
  assign tmp727 = (tmp484 & tmp605) | (tmp484 & tmp726) | (tmp605 & tmp726);
  wire tmp728;
  assign tmp728 = 1'b0;
  wire tmp729;
  assign tmp729 = 1'b0;
  wire tmp730;
  assign tmp730 = 1'b0;
  wire tmp731;
  assign tmp731 = (tmp728 & tmp729) | (tmp728 & tmp730) | (tmp729 & tmp730);
  wire tmp732;
  assign tmp732 = 1'b0;
  wire tmp733;
  assign tmp733 = 1'b0;
  wire tmp734;
  assign tmp734 = 1'b0;
  wire tmp735;
  assign tmp735 = (tmp732 & tmp733) | (tmp732 & tmp734) | (tmp733 & tmp734);
  wire tmp736;
  assign tmp736 = 1'b0;
  wire tmp737;
  assign tmp737 = 1'b0;
  wire tmp738;
  assign tmp738 = 1'b0;
  wire tmp739;
  assign tmp739 = (tmp736 & tmp737) | (tmp736 & tmp738) | (tmp737 & tmp738);
  wire tmp740;
  assign tmp740 = (tmp731 & tmp735) | (tmp731 & tmp739) | (tmp735 & tmp739);
  wire tmp741;
  assign tmp741 = 1'b0;
  wire tmp742;
  assign tmp742 = 1'b0;
  wire tmp743;
  assign tmp743 = 1'b0;
  wire tmp744;
  assign tmp744 = (tmp741 & tmp742) | (tmp741 & tmp743) | (tmp742 & tmp743);
  wire tmp745;
  assign tmp745 = 1'b0;
  wire tmp746;
  assign tmp746 = 1'b0;
  wire tmp747;
  assign tmp747 = 1'b0;
  wire tmp748;
  assign tmp748 = (tmp745 & tmp746) | (tmp745 & tmp747) | (tmp746 & tmp747);
  wire tmp749;
  assign tmp749 = 1'b0;
  wire tmp750;
  assign tmp750 = 1'b0;
  wire tmp751;
  assign tmp751 = 1'b0;
  wire tmp752;
  assign tmp752 = (tmp749 & tmp750) | (tmp749 & tmp751) | (tmp750 & tmp751);
  wire tmp753;
  assign tmp753 = (tmp744 & tmp748) | (tmp744 & tmp752) | (tmp748 & tmp752);
  wire tmp754;
  assign tmp754 = 1'b0;
  wire tmp755;
  assign tmp755 = 1'b0;
  wire tmp756;
  assign tmp756 = 1'b0;
  wire tmp757;
  assign tmp757 = (tmp754 & tmp755) | (tmp754 & tmp756) | (tmp755 & tmp756);
  wire tmp758;
  assign tmp758 = 1'b0;
  wire tmp759;
  assign tmp759 = 1'b0;
  wire tmp760;
  assign tmp760 = 1'b0;
  wire tmp761;
  assign tmp761 = (tmp758 & tmp759) | (tmp758 & tmp760) | (tmp759 & tmp760);
  wire tmp762;
  assign tmp762 = 1'b0;
  wire tmp763;
  assign tmp763 = 1'b0;
  wire tmp764;
  assign tmp764 = 1'b0;
  wire tmp765;
  assign tmp765 = (tmp762 & tmp763) | (tmp762 & tmp764) | (tmp763 & tmp764);
  wire tmp766;
  assign tmp766 = (tmp757 & tmp761) | (tmp757 & tmp765) | (tmp761 & tmp765);
  wire tmp767;
  assign tmp767 = (tmp740 & tmp753) | (tmp740 & tmp766) | (tmp753 & tmp766);
  wire tmp768;
  assign tmp768 = 1'b0;
  wire tmp769;
  assign tmp769 = 1'b0;
  wire tmp770;
  assign tmp770 = 1'b0;
  wire tmp771;
  assign tmp771 = (tmp768 & tmp769) | (tmp768 & tmp770) | (tmp769 & tmp770);
  wire tmp772;
  assign tmp772 = 1'b0;
  wire tmp773;
  assign tmp773 = 1'b0;
  wire tmp774;
  assign tmp774 = 1'b0;
  wire tmp775;
  assign tmp775 = (tmp772 & tmp773) | (tmp772 & tmp774) | (tmp773 & tmp774);
  wire tmp776;
  assign tmp776 = 1'b0;
  wire tmp777;
  assign tmp777 = 1'b0;
  wire tmp778;
  assign tmp778 = 1'b0;
  wire tmp779;
  assign tmp779 = (tmp776 & tmp777) | (tmp776 & tmp778) | (tmp777 & tmp778);
  wire tmp780;
  assign tmp780 = (tmp771 & tmp775) | (tmp771 & tmp779) | (tmp775 & tmp779);
  wire tmp781;
  assign tmp781 = 1'b0;
  wire tmp782;
  assign tmp782 = 1'b0;
  wire tmp783;
  assign tmp783 = 1'b0;
  wire tmp784;
  assign tmp784 = (tmp781 & tmp782) | (tmp781 & tmp783) | (tmp782 & tmp783);
  wire tmp785;
  assign tmp785 = 1'b0;
  wire tmp786;
  assign tmp786 = 1'b1;
  wire tmp787;
  assign tmp787 = 1'b0;
  wire tmp788;
  assign tmp788 = (tmp785 & tmp786) | (tmp785 & tmp787) | (tmp786 & tmp787);
  wire tmp789;
  assign tmp789 = 1'b0;
  wire tmp790;
  assign tmp790 = 1'b0;
  wire tmp791;
  assign tmp791 = 1'b0;
  wire tmp792;
  assign tmp792 = (tmp789 & tmp790) | (tmp789 & tmp791) | (tmp790 & tmp791);
  wire tmp793;
  assign tmp793 = (tmp784 & tmp788) | (tmp784 & tmp792) | (tmp788 & tmp792);
  wire tmp794;
  assign tmp794 = 1'b0;
  wire tmp795;
  assign tmp795 = 1'b0;
  wire tmp796;
  assign tmp796 = 1'b0;
  wire tmp797;
  assign tmp797 = (tmp794 & tmp795) | (tmp794 & tmp796) | (tmp795 & tmp796);
  wire tmp798;
  assign tmp798 = 1'b0;
  wire tmp799;
  assign tmp799 = 1'b0;
  wire tmp800;
  assign tmp800 = 1'b0;
  wire tmp801;
  assign tmp801 = (tmp798 & tmp799) | (tmp798 & tmp800) | (tmp799 & tmp800);
  wire tmp802;
  assign tmp802 = 1'b0;
  wire tmp803;
  assign tmp803 = 1'b0;
  wire tmp804;
  assign tmp804 = 1'b0;
  wire tmp805;
  assign tmp805 = (tmp802 & tmp803) | (tmp802 & tmp804) | (tmp803 & tmp804);
  wire tmp806;
  assign tmp806 = (tmp797 & tmp801) | (tmp797 & tmp805) | (tmp801 & tmp805);
  wire tmp807;
  assign tmp807 = (tmp780 & tmp793) | (tmp780 & tmp806) | (tmp793 & tmp806);
  wire tmp808;
  assign tmp808 = 1'b0;
  wire tmp809;
  assign tmp809 = 1'b0;
  wire tmp810;
  assign tmp810 = 1'b0;
  wire tmp811;
  assign tmp811 = (tmp808 & tmp809) | (tmp808 & tmp810) | (tmp809 & tmp810);
  wire tmp812;
  assign tmp812 = 1'b0;
  wire tmp813;
  assign tmp813 = 1'b0;
  wire tmp814;
  assign tmp814 = 1'b0;
  wire tmp815;
  assign tmp815 = (tmp812 & tmp813) | (tmp812 & tmp814) | (tmp813 & tmp814);
  wire tmp816;
  assign tmp816 = 1'b0;
  wire tmp817;
  assign tmp817 = 1'b0;
  wire tmp818;
  assign tmp818 = 1'b0;
  wire tmp819;
  assign tmp819 = (tmp816 & tmp817) | (tmp816 & tmp818) | (tmp817 & tmp818);
  wire tmp820;
  assign tmp820 = (tmp811 & tmp815) | (tmp811 & tmp819) | (tmp815 & tmp819);
  wire tmp821;
  assign tmp821 = 1'b0;
  wire tmp822;
  assign tmp822 = 1'b0;
  wire tmp823;
  assign tmp823 = 1'b0;
  wire tmp824;
  assign tmp824 = (tmp821 & tmp822) | (tmp821 & tmp823) | (tmp822 & tmp823);
  wire tmp825;
  assign tmp825 = 1'b0;
  wire tmp826;
  assign tmp826 = 1'b0;
  wire tmp827;
  assign tmp827 = 1'b0;
  wire tmp828;
  assign tmp828 = (tmp825 & tmp826) | (tmp825 & tmp827) | (tmp826 & tmp827);
  wire tmp829;
  assign tmp829 = 1'b0;
  wire tmp830;
  assign tmp830 = 1'b0;
  wire tmp831;
  assign tmp831 = 1'b0;
  wire tmp832;
  assign tmp832 = (tmp829 & tmp830) | (tmp829 & tmp831) | (tmp830 & tmp831);
  wire tmp833;
  assign tmp833 = (tmp824 & tmp828) | (tmp824 & tmp832) | (tmp828 & tmp832);
  wire tmp834;
  assign tmp834 = 1'b0;
  wire tmp835;
  assign tmp835 = 1'b0;
  wire tmp836;
  assign tmp836 = 1'b0;
  wire tmp837;
  assign tmp837 = (tmp834 & tmp835) | (tmp834 & tmp836) | (tmp835 & tmp836);
  wire tmp838;
  assign tmp838 = 1'b0;
  wire tmp839;
  assign tmp839 = 1'b0;
  wire tmp840;
  assign tmp840 = 1'b0;
  wire tmp841;
  assign tmp841 = (tmp838 & tmp839) | (tmp838 & tmp840) | (tmp839 & tmp840);
  wire tmp842;
  assign tmp842 = 1'b0;
  wire tmp843;
  assign tmp843 = 1'b0;
  wire tmp844;
  assign tmp844 = 1'b0;
  wire tmp845;
  assign tmp845 = (tmp842 & tmp843) | (tmp842 & tmp844) | (tmp843 & tmp844);
  wire tmp846;
  assign tmp846 = (tmp837 & tmp841) | (tmp837 & tmp845) | (tmp841 & tmp845);
  wire tmp847;
  assign tmp847 = (tmp820 & tmp833) | (tmp820 & tmp846) | (tmp833 & tmp846);
  wire tmp848;
  assign tmp848 = (tmp767 & tmp807) | (tmp767 & tmp847) | (tmp807 & tmp847);
  wire tmp849;
  assign tmp849 = 1'b0;
  wire tmp850;
  assign tmp850 = 1'b0;
  wire tmp851;
  assign tmp851 = 1'b0;
  wire tmp852;
  assign tmp852 = (tmp849 & tmp850) | (tmp849 & tmp851) | (tmp850 & tmp851);
  wire tmp853;
  assign tmp853 = 1'b0;
  wire tmp854;
  assign tmp854 = 1'b0;
  wire tmp855;
  assign tmp855 = 1'b0;
  wire tmp856;
  assign tmp856 = (tmp853 & tmp854) | (tmp853 & tmp855) | (tmp854 & tmp855);
  wire tmp857;
  assign tmp857 = 1'b0;
  wire tmp858;
  assign tmp858 = 1'b0;
  wire tmp859;
  assign tmp859 = 1'b0;
  wire tmp860;
  assign tmp860 = (tmp857 & tmp858) | (tmp857 & tmp859) | (tmp858 & tmp859);
  wire tmp861;
  assign tmp861 = (tmp852 & tmp856) | (tmp852 & tmp860) | (tmp856 & tmp860);
  wire tmp862;
  assign tmp862 = 1'b0;
  wire tmp863;
  assign tmp863 = 1'b0;
  wire tmp864;
  assign tmp864 = 1'b0;
  wire tmp865;
  assign tmp865 = (tmp862 & tmp863) | (tmp862 & tmp864) | (tmp863 & tmp864);
  wire tmp866;
  assign tmp866 = 1'b0;
  wire tmp867;
  assign tmp867 = 1'b1;
  wire tmp868;
  assign tmp868 = 1'b0;
  wire tmp869;
  assign tmp869 = (tmp866 & tmp867) | (tmp866 & tmp868) | (tmp867 & tmp868);
  wire tmp870;
  assign tmp870 = 1'b0;
  wire tmp871;
  assign tmp871 = 1'b0;
  wire tmp872;
  assign tmp872 = 1'b0;
  wire tmp873;
  assign tmp873 = (tmp870 & tmp871) | (tmp870 & tmp872) | (tmp871 & tmp872);
  wire tmp874;
  assign tmp874 = (tmp865 & tmp869) | (tmp865 & tmp873) | (tmp869 & tmp873);
  wire tmp875;
  assign tmp875 = 1'b0;
  wire tmp876;
  assign tmp876 = 1'b0;
  wire tmp877;
  assign tmp877 = 1'b0;
  wire tmp878;
  assign tmp878 = (tmp875 & tmp876) | (tmp875 & tmp877) | (tmp876 & tmp877);
  wire tmp879;
  assign tmp879 = 1'b0;
  wire tmp880;
  assign tmp880 = 1'b0;
  wire tmp881;
  assign tmp881 = 1'b0;
  wire tmp882;
  assign tmp882 = (tmp879 & tmp880) | (tmp879 & tmp881) | (tmp880 & tmp881);
  wire tmp883;
  assign tmp883 = 1'b0;
  wire tmp884;
  assign tmp884 = 1'b0;
  wire tmp885;
  assign tmp885 = 1'b0;
  wire tmp886;
  assign tmp886 = (tmp883 & tmp884) | (tmp883 & tmp885) | (tmp884 & tmp885);
  wire tmp887;
  assign tmp887 = (tmp878 & tmp882) | (tmp878 & tmp886) | (tmp882 & tmp886);
  wire tmp888;
  assign tmp888 = (tmp861 & tmp874) | (tmp861 & tmp887) | (tmp874 & tmp887);
  wire tmp889;
  assign tmp889 = 1'b0;
  wire tmp890;
  assign tmp890 = 1'b0;
  wire tmp891;
  assign tmp891 = 1'b0;
  wire tmp892;
  assign tmp892 = (tmp889 & tmp890) | (tmp889 & tmp891) | (tmp890 & tmp891);
  wire tmp893;
  assign tmp893 = 1'b0;
  wire tmp894;
  assign tmp894 = 1'b1;
  wire tmp895;
  assign tmp895 = 1'b0;
  wire tmp896;
  assign tmp896 = (tmp893 & tmp894) | (tmp893 & tmp895) | (tmp894 & tmp895);
  wire tmp897;
  assign tmp897 = 1'b0;
  wire tmp898;
  assign tmp898 = 1'b0;
  wire tmp899;
  assign tmp899 = 1'b0;
  wire tmp900;
  assign tmp900 = (tmp897 & tmp898) | (tmp897 & tmp899) | (tmp898 & tmp899);
  wire tmp901;
  assign tmp901 = (tmp892 & tmp896) | (tmp892 & tmp900) | (tmp896 & tmp900);
  wire tmp902;
  assign tmp902 = 1'b0;
  wire tmp903;
  assign tmp903 = 1'b1;
  wire tmp904;
  assign tmp904 = 1'b0;
  wire tmp905;
  assign tmp905 = (tmp902 & tmp903) | (tmp902 & tmp904) | (tmp903 & tmp904);
  wire tmp906;
  assign tmp906 = 1'b1;
  wire tmp907;
  assign tmp907 = 1'b1;
  wire tmp908;
  assign tmp908 = 1'b1;
  wire tmp909;
  assign tmp909 = (tmp906 & tmp907) | (tmp906 & tmp908) | (tmp907 & tmp908);
  wire tmp910;
  assign tmp910 = 1'b0;
  wire tmp911;
  assign tmp911 = 1'b1;
  wire tmp912;
  assign tmp912 = 1'b0;
  wire tmp913;
  assign tmp913 = (tmp910 & tmp911) | (tmp910 & tmp912) | (tmp911 & tmp912);
  wire tmp914;
  assign tmp914 = (tmp905 & tmp909) | (tmp905 & tmp913) | (tmp909 & tmp913);
  wire tmp915;
  assign tmp915 = 1'b0;
  wire tmp916;
  assign tmp916 = 1'b0;
  wire tmp917;
  assign tmp917 = 1'b0;
  wire tmp918;
  assign tmp918 = (tmp915 & tmp916) | (tmp915 & tmp917) | (tmp916 & tmp917);
  wire tmp919;
  assign tmp919 = 1'b0;
  wire tmp920;
  assign tmp920 = 1'b1;
  wire tmp921;
  assign tmp921 = 1'b0;
  wire tmp922;
  assign tmp922 = (tmp919 & tmp920) | (tmp919 & tmp921) | (tmp920 & tmp921);
  wire tmp923;
  assign tmp923 = 1'b0;
  wire tmp924;
  assign tmp924 = 1'b0;
  wire tmp925;
  assign tmp925 = 1'b0;
  wire tmp926;
  assign tmp926 = (tmp923 & tmp924) | (tmp923 & tmp925) | (tmp924 & tmp925);
  wire tmp927;
  assign tmp927 = (tmp918 & tmp922) | (tmp918 & tmp926) | (tmp922 & tmp926);
  wire tmp928;
  assign tmp928 = (tmp901 & tmp914) | (tmp901 & tmp927) | (tmp914 & tmp927);
  wire tmp929;
  assign tmp929 = 1'b0;
  wire tmp930;
  assign tmp930 = 1'b0;
  wire tmp931;
  assign tmp931 = 1'b0;
  wire tmp932;
  assign tmp932 = (tmp929 & tmp930) | (tmp929 & tmp931) | (tmp930 & tmp931);
  wire tmp933;
  assign tmp933 = 1'b0;
  wire tmp934;
  assign tmp934 = 1'b0;
  wire tmp935;
  assign tmp935 = 1'b0;
  wire tmp936;
  assign tmp936 = (tmp933 & tmp934) | (tmp933 & tmp935) | (tmp934 & tmp935);
  wire tmp937;
  assign tmp937 = 1'b0;
  wire tmp938;
  assign tmp938 = 1'b0;
  wire tmp939;
  assign tmp939 = 1'b0;
  wire tmp940;
  assign tmp940 = (tmp937 & tmp938) | (tmp937 & tmp939) | (tmp938 & tmp939);
  wire tmp941;
  assign tmp941 = (tmp932 & tmp936) | (tmp932 & tmp940) | (tmp936 & tmp940);
  wire tmp942;
  assign tmp942 = 1'b0;
  wire tmp943;
  assign tmp943 = 1'b0;
  wire tmp944;
  assign tmp944 = 1'b0;
  wire tmp945;
  assign tmp945 = (tmp942 & tmp943) | (tmp942 & tmp944) | (tmp943 & tmp944);
  wire tmp946;
  assign tmp946 = 1'b0;
  wire tmp947;
  assign tmp947 = 1'b1;
  wire tmp948;
  assign tmp948 = 1'b0;
  wire tmp949;
  assign tmp949 = (tmp946 & tmp947) | (tmp946 & tmp948) | (tmp947 & tmp948);
  wire tmp950;
  assign tmp950 = 1'b0;
  wire tmp951;
  assign tmp951 = 1'b0;
  wire tmp952;
  assign tmp952 = 1'b0;
  wire tmp953;
  assign tmp953 = (tmp950 & tmp951) | (tmp950 & tmp952) | (tmp951 & tmp952);
  wire tmp954;
  assign tmp954 = (tmp945 & tmp949) | (tmp945 & tmp953) | (tmp949 & tmp953);
  wire tmp955;
  assign tmp955 = 1'b0;
  wire tmp956;
  assign tmp956 = 1'b0;
  wire tmp957;
  assign tmp957 = 1'b0;
  wire tmp958;
  assign tmp958 = (tmp955 & tmp956) | (tmp955 & tmp957) | (tmp956 & tmp957);
  wire tmp959;
  assign tmp959 = 1'b0;
  wire tmp960;
  assign tmp960 = 1'b0;
  wire tmp961;
  assign tmp961 = 1'b0;
  wire tmp962;
  assign tmp962 = (tmp959 & tmp960) | (tmp959 & tmp961) | (tmp960 & tmp961);
  wire tmp963;
  assign tmp963 = 1'b0;
  wire tmp964;
  assign tmp964 = 1'b0;
  wire tmp965;
  assign tmp965 = 1'b0;
  wire tmp966;
  assign tmp966 = (tmp963 & tmp964) | (tmp963 & tmp965) | (tmp964 & tmp965);
  wire tmp967;
  assign tmp967 = (tmp958 & tmp962) | (tmp958 & tmp966) | (tmp962 & tmp966);
  wire tmp968;
  assign tmp968 = (tmp941 & tmp954) | (tmp941 & tmp967) | (tmp954 & tmp967);
  wire tmp969;
  assign tmp969 = (tmp888 & tmp928) | (tmp888 & tmp968) | (tmp928 & tmp968);
  wire tmp970;
  assign tmp970 = 1'b0;
  wire tmp971;
  assign tmp971 = 1'b0;
  wire tmp972;
  assign tmp972 = 1'b0;
  wire tmp973;
  assign tmp973 = (tmp970 & tmp971) | (tmp970 & tmp972) | (tmp971 & tmp972);
  wire tmp974;
  assign tmp974 = 1'b0;
  wire tmp975;
  assign tmp975 = 1'b0;
  wire tmp976;
  assign tmp976 = 1'b0;
  wire tmp977;
  assign tmp977 = (tmp974 & tmp975) | (tmp974 & tmp976) | (tmp975 & tmp976);
  wire tmp978;
  assign tmp978 = 1'b0;
  wire tmp979;
  assign tmp979 = 1'b0;
  wire tmp980;
  assign tmp980 = 1'b0;
  wire tmp981;
  assign tmp981 = (tmp978 & tmp979) | (tmp978 & tmp980) | (tmp979 & tmp980);
  wire tmp982;
  assign tmp982 = (tmp973 & tmp977) | (tmp973 & tmp981) | (tmp977 & tmp981);
  wire tmp983;
  assign tmp983 = 1'b0;
  wire tmp984;
  assign tmp984 = 1'b0;
  wire tmp985;
  assign tmp985 = 1'b0;
  wire tmp986;
  assign tmp986 = (tmp983 & tmp984) | (tmp983 & tmp985) | (tmp984 & tmp985);
  wire tmp987;
  assign tmp987 = 1'b0;
  wire tmp988;
  assign tmp988 = 1'b0;
  wire tmp989;
  assign tmp989 = 1'b0;
  wire tmp990;
  assign tmp990 = (tmp987 & tmp988) | (tmp987 & tmp989) | (tmp988 & tmp989);
  wire tmp991;
  assign tmp991 = 1'b0;
  wire tmp992;
  assign tmp992 = 1'b0;
  wire tmp993;
  assign tmp993 = 1'b0;
  wire tmp994;
  assign tmp994 = (tmp991 & tmp992) | (tmp991 & tmp993) | (tmp992 & tmp993);
  wire tmp995;
  assign tmp995 = (tmp986 & tmp990) | (tmp986 & tmp994) | (tmp990 & tmp994);
  wire tmp996;
  assign tmp996 = 1'b0;
  wire tmp997;
  assign tmp997 = 1'b0;
  wire tmp998;
  assign tmp998 = 1'b0;
  wire tmp999;
  assign tmp999 = (tmp996 & tmp997) | (tmp996 & tmp998) | (tmp997 & tmp998);
  wire tmp1000;
  assign tmp1000 = 1'b0;
  wire tmp1001;
  assign tmp1001 = 1'b0;
  wire tmp1002;
  assign tmp1002 = 1'b0;
  wire tmp1003;
  assign tmp1003 = (tmp1000 & tmp1001) | (tmp1000 & tmp1002) | (tmp1001 & tmp1002);
  wire tmp1004;
  assign tmp1004 = 1'b0;
  wire tmp1005;
  assign tmp1005 = 1'b0;
  wire tmp1006;
  assign tmp1006 = 1'b0;
  wire tmp1007;
  assign tmp1007 = (tmp1004 & tmp1005) | (tmp1004 & tmp1006) | (tmp1005 & tmp1006);
  wire tmp1008;
  assign tmp1008 = (tmp999 & tmp1003) | (tmp999 & tmp1007) | (tmp1003 & tmp1007);
  wire tmp1009;
  assign tmp1009 = (tmp982 & tmp995) | (tmp982 & tmp1008) | (tmp995 & tmp1008);
  wire tmp1010;
  assign tmp1010 = 1'b0;
  wire tmp1011;
  assign tmp1011 = 1'b0;
  wire tmp1012;
  assign tmp1012 = 1'b0;
  wire tmp1013;
  assign tmp1013 = (tmp1010 & tmp1011) | (tmp1010 & tmp1012) | (tmp1011 & tmp1012);
  wire tmp1014;
  assign tmp1014 = 1'b0;
  wire tmp1015;
  assign tmp1015 = 1'b0;
  wire tmp1016;
  assign tmp1016 = 1'b0;
  wire tmp1017;
  assign tmp1017 = (tmp1014 & tmp1015) | (tmp1014 & tmp1016) | (tmp1015 & tmp1016);
  wire tmp1018;
  assign tmp1018 = 1'b0;
  wire tmp1019;
  assign tmp1019 = 1'b0;
  wire tmp1020;
  assign tmp1020 = 1'b0;
  wire tmp1021;
  assign tmp1021 = (tmp1018 & tmp1019) | (tmp1018 & tmp1020) | (tmp1019 & tmp1020);
  wire tmp1022;
  assign tmp1022 = (tmp1013 & tmp1017) | (tmp1013 & tmp1021) | (tmp1017 & tmp1021);
  wire tmp1023;
  assign tmp1023 = 1'b0;
  wire tmp1024;
  assign tmp1024 = 1'b0;
  wire tmp1025;
  assign tmp1025 = 1'b0;
  wire tmp1026;
  assign tmp1026 = (tmp1023 & tmp1024) | (tmp1023 & tmp1025) | (tmp1024 & tmp1025);
  wire tmp1027;
  assign tmp1027 = 1'b0;
  wire tmp1028;
  assign tmp1028 = 1'b1;
  wire tmp1029;
  assign tmp1029 = 1'b0;
  wire tmp1030;
  assign tmp1030 = (tmp1027 & tmp1028) | (tmp1027 & tmp1029) | (tmp1028 & tmp1029);
  wire tmp1031;
  assign tmp1031 = 1'b0;
  wire tmp1032;
  assign tmp1032 = 1'b0;
  wire tmp1033;
  assign tmp1033 = 1'b0;
  wire tmp1034;
  assign tmp1034 = (tmp1031 & tmp1032) | (tmp1031 & tmp1033) | (tmp1032 & tmp1033);
  wire tmp1035;
  assign tmp1035 = (tmp1026 & tmp1030) | (tmp1026 & tmp1034) | (tmp1030 & tmp1034);
  wire tmp1036;
  assign tmp1036 = 1'b0;
  wire tmp1037;
  assign tmp1037 = 1'b0;
  wire tmp1038;
  assign tmp1038 = 1'b0;
  wire tmp1039;
  assign tmp1039 = (tmp1036 & tmp1037) | (tmp1036 & tmp1038) | (tmp1037 & tmp1038);
  wire tmp1040;
  assign tmp1040 = 1'b0;
  wire tmp1041;
  assign tmp1041 = 1'b0;
  wire tmp1042;
  assign tmp1042 = 1'b0;
  wire tmp1043;
  assign tmp1043 = (tmp1040 & tmp1041) | (tmp1040 & tmp1042) | (tmp1041 & tmp1042);
  wire tmp1044;
  assign tmp1044 = 1'b0;
  wire tmp1045;
  assign tmp1045 = 1'b0;
  wire tmp1046;
  assign tmp1046 = 1'b0;
  wire tmp1047;
  assign tmp1047 = (tmp1044 & tmp1045) | (tmp1044 & tmp1046) | (tmp1045 & tmp1046);
  wire tmp1048;
  assign tmp1048 = (tmp1039 & tmp1043) | (tmp1039 & tmp1047) | (tmp1043 & tmp1047);
  wire tmp1049;
  assign tmp1049 = (tmp1022 & tmp1035) | (tmp1022 & tmp1048) | (tmp1035 & tmp1048);
  wire tmp1050;
  assign tmp1050 = 1'b0;
  wire tmp1051;
  assign tmp1051 = 1'b0;
  wire tmp1052;
  assign tmp1052 = 1'b0;
  wire tmp1053;
  assign tmp1053 = (tmp1050 & tmp1051) | (tmp1050 & tmp1052) | (tmp1051 & tmp1052);
  wire tmp1054;
  assign tmp1054 = 1'b0;
  wire tmp1055;
  assign tmp1055 = 1'b0;
  wire tmp1056;
  assign tmp1056 = 1'b0;
  wire tmp1057;
  assign tmp1057 = (tmp1054 & tmp1055) | (tmp1054 & tmp1056) | (tmp1055 & tmp1056);
  wire tmp1058;
  assign tmp1058 = 1'b0;
  wire tmp1059;
  assign tmp1059 = 1'b0;
  wire tmp1060;
  assign tmp1060 = 1'b0;
  wire tmp1061;
  assign tmp1061 = (tmp1058 & tmp1059) | (tmp1058 & tmp1060) | (tmp1059 & tmp1060);
  wire tmp1062;
  assign tmp1062 = (tmp1053 & tmp1057) | (tmp1053 & tmp1061) | (tmp1057 & tmp1061);
  wire tmp1063;
  assign tmp1063 = 1'b0;
  wire tmp1064;
  assign tmp1064 = 1'b0;
  wire tmp1065;
  assign tmp1065 = 1'b0;
  wire tmp1066;
  assign tmp1066 = (tmp1063 & tmp1064) | (tmp1063 & tmp1065) | (tmp1064 & tmp1065);
  wire tmp1067;
  assign tmp1067 = 1'b0;
  wire tmp1068;
  assign tmp1068 = 1'b0;
  wire tmp1069;
  assign tmp1069 = 1'b0;
  wire tmp1070;
  assign tmp1070 = (tmp1067 & tmp1068) | (tmp1067 & tmp1069) | (tmp1068 & tmp1069);
  wire tmp1071;
  assign tmp1071 = 1'b0;
  wire tmp1072;
  assign tmp1072 = 1'b0;
  wire tmp1073;
  assign tmp1073 = 1'b0;
  wire tmp1074;
  assign tmp1074 = (tmp1071 & tmp1072) | (tmp1071 & tmp1073) | (tmp1072 & tmp1073);
  wire tmp1075;
  assign tmp1075 = (tmp1066 & tmp1070) | (tmp1066 & tmp1074) | (tmp1070 & tmp1074);
  wire tmp1076;
  assign tmp1076 = 1'b0;
  wire tmp1077;
  assign tmp1077 = 1'b0;
  wire tmp1078;
  assign tmp1078 = 1'b0;
  wire tmp1079;
  assign tmp1079 = (tmp1076 & tmp1077) | (tmp1076 & tmp1078) | (tmp1077 & tmp1078);
  wire tmp1080;
  assign tmp1080 = 1'b0;
  wire tmp1081;
  assign tmp1081 = 1'b0;
  wire tmp1082;
  assign tmp1082 = 1'b0;
  wire tmp1083;
  assign tmp1083 = (tmp1080 & tmp1081) | (tmp1080 & tmp1082) | (tmp1081 & tmp1082);
  wire tmp1084;
  assign tmp1084 = 1'b0;
  wire tmp1085;
  assign tmp1085 = 1'b0;
  wire tmp1086;
  assign tmp1086 = 1'b0;
  wire tmp1087;
  assign tmp1087 = (tmp1084 & tmp1085) | (tmp1084 & tmp1086) | (tmp1085 & tmp1086);
  wire tmp1088;
  assign tmp1088 = (tmp1079 & tmp1083) | (tmp1079 & tmp1087) | (tmp1083 & tmp1087);
  wire tmp1089;
  assign tmp1089 = (tmp1062 & tmp1075) | (tmp1062 & tmp1088) | (tmp1075 & tmp1088);
  wire tmp1090;
  assign tmp1090 = (tmp1009 & tmp1049) | (tmp1009 & tmp1089) | (tmp1049 & tmp1089);
  wire tmp1091;
  assign tmp1091 = (tmp848 & tmp969) | (tmp848 & tmp1090) | (tmp969 & tmp1090);
  wire tmp1092;
  assign tmp1092 = (tmp363 & tmp727) | (tmp363 & tmp1091) | (tmp727 & tmp1091);
  wire tmp1093;
  assign tmp1093 = pi1;
  wire tmp1094;
  assign tmp1094 = pi2;
  wire tmp1095;
  assign tmp1095 = 1'b0;
  wire tmp1096;
  assign tmp1096 = (tmp1093 & tmp1094) | (tmp1093 & tmp1095) | (tmp1094 & tmp1095);
  wire tmp1097;
  assign tmp1097 = pi2;
  wire tmp1098;
  assign tmp1098 = pi3;
  wire tmp1099;
  assign tmp1099 = 1'b0;
  wire tmp1100;
  assign tmp1100 = (tmp1097 & tmp1098) | (tmp1097 & tmp1099) | (tmp1098 & tmp1099);
  wire tmp1101;
  assign tmp1101 = 1'b0;
  wire tmp1102;
  assign tmp1102 = 1'b0;
  wire tmp1103;
  assign tmp1103 = 1'b0;
  wire tmp1104;
  assign tmp1104 = (tmp1101 & tmp1102) | (tmp1101 & tmp1103) | (tmp1102 & tmp1103);
  wire tmp1105;
  assign tmp1105 = (tmp1096 & tmp1100) | (tmp1096 & tmp1104) | (tmp1100 & tmp1104);
  wire tmp1106;
  assign tmp1106 = pi2;
  wire tmp1107;
  assign tmp1107 = pi3;
  wire tmp1108;
  assign tmp1108 = 1'b0;
  wire tmp1109;
  assign tmp1109 = (tmp1106 & tmp1107) | (tmp1106 & tmp1108) | (tmp1107 & tmp1108);
  wire tmp1110;
  assign tmp1110 = pi3;
  wire tmp1111;
  assign tmp1111 = 1'b1;
  wire tmp1112;
  assign tmp1112 = 1'b0;
  wire tmp1113;
  assign tmp1113 = (tmp1110 & tmp1111) | (tmp1110 & tmp1112) | (tmp1111 & tmp1112);
  wire tmp1114;
  assign tmp1114 = 1'b0;
  wire tmp1115;
  assign tmp1115 = 1'b0;
  wire tmp1116;
  assign tmp1116 = 1'b0;
  wire tmp1117;
  assign tmp1117 = (tmp1114 & tmp1115) | (tmp1114 & tmp1116) | (tmp1115 & tmp1116);
  wire tmp1118;
  assign tmp1118 = (tmp1109 & tmp1113) | (tmp1109 & tmp1117) | (tmp1113 & tmp1117);
  wire tmp1119;
  assign tmp1119 = 1'b0;
  wire tmp1120;
  assign tmp1120 = 1'b0;
  wire tmp1121;
  assign tmp1121 = 1'b0;
  wire tmp1122;
  assign tmp1122 = (tmp1119 & tmp1120) | (tmp1119 & tmp1121) | (tmp1120 & tmp1121);
  wire tmp1123;
  assign tmp1123 = 1'b0;
  wire tmp1124;
  assign tmp1124 = 1'b0;
  wire tmp1125;
  assign tmp1125 = 1'b0;
  wire tmp1126;
  assign tmp1126 = (tmp1123 & tmp1124) | (tmp1123 & tmp1125) | (tmp1124 & tmp1125);
  wire tmp1127;
  assign tmp1127 = 1'b0;
  wire tmp1128;
  assign tmp1128 = 1'b0;
  wire tmp1129;
  assign tmp1129 = 1'b0;
  wire tmp1130;
  assign tmp1130 = (tmp1127 & tmp1128) | (tmp1127 & tmp1129) | (tmp1128 & tmp1129);
  wire tmp1131;
  assign tmp1131 = (tmp1122 & tmp1126) | (tmp1122 & tmp1130) | (tmp1126 & tmp1130);
  wire tmp1132;
  assign tmp1132 = (tmp1105 & tmp1118) | (tmp1105 & tmp1131) | (tmp1118 & tmp1131);
  wire tmp1133;
  assign tmp1133 = pi2;
  wire tmp1134;
  assign tmp1134 = pi3;
  wire tmp1135;
  assign tmp1135 = 1'b0;
  wire tmp1136;
  assign tmp1136 = (tmp1133 & tmp1134) | (tmp1133 & tmp1135) | (tmp1134 & tmp1135);
  wire tmp1137;
  assign tmp1137 = pi3;
  wire tmp1138;
  assign tmp1138 = 1'b1;
  wire tmp1139;
  assign tmp1139 = 1'b0;
  wire tmp1140;
  assign tmp1140 = (tmp1137 & tmp1138) | (tmp1137 & tmp1139) | (tmp1138 & tmp1139);
  wire tmp1141;
  assign tmp1141 = 1'b0;
  wire tmp1142;
  assign tmp1142 = 1'b0;
  wire tmp1143;
  assign tmp1143 = 1'b0;
  wire tmp1144;
  assign tmp1144 = (tmp1141 & tmp1142) | (tmp1141 & tmp1143) | (tmp1142 & tmp1143);
  wire tmp1145;
  assign tmp1145 = (tmp1136 & tmp1140) | (tmp1136 & tmp1144) | (tmp1140 & tmp1144);
  wire tmp1146;
  assign tmp1146 = pi3;
  wire tmp1147;
  assign tmp1147 = 1'b1;
  wire tmp1148;
  assign tmp1148 = 1'b0;
  wire tmp1149;
  assign tmp1149 = (tmp1146 & tmp1147) | (tmp1146 & tmp1148) | (tmp1147 & tmp1148);
  wire tmp1150;
  assign tmp1150 = 1'b1;
  wire tmp1151;
  assign tmp1151 = 1'b1;
  wire tmp1152;
  assign tmp1152 = 1'b1;
  wire tmp1153;
  assign tmp1153 = (tmp1150 & tmp1151) | (tmp1150 & tmp1152) | (tmp1151 & tmp1152);
  wire tmp1154;
  assign tmp1154 = 1'b0;
  wire tmp1155;
  assign tmp1155 = 1'b1;
  wire tmp1156;
  assign tmp1156 = 1'b0;
  wire tmp1157;
  assign tmp1157 = (tmp1154 & tmp1155) | (tmp1154 & tmp1156) | (tmp1155 & tmp1156);
  wire tmp1158;
  assign tmp1158 = (tmp1149 & tmp1153) | (tmp1149 & tmp1157) | (tmp1153 & tmp1157);
  wire tmp1159;
  assign tmp1159 = 1'b0;
  wire tmp1160;
  assign tmp1160 = 1'b0;
  wire tmp1161;
  assign tmp1161 = 1'b0;
  wire tmp1162;
  assign tmp1162 = (tmp1159 & tmp1160) | (tmp1159 & tmp1161) | (tmp1160 & tmp1161);
  wire tmp1163;
  assign tmp1163 = 1'b0;
  wire tmp1164;
  assign tmp1164 = 1'b1;
  wire tmp1165;
  assign tmp1165 = 1'b0;
  wire tmp1166;
  assign tmp1166 = (tmp1163 & tmp1164) | (tmp1163 & tmp1165) | (tmp1164 & tmp1165);
  wire tmp1167;
  assign tmp1167 = 1'b0;
  wire tmp1168;
  assign tmp1168 = 1'b0;
  wire tmp1169;
  assign tmp1169 = 1'b0;
  wire tmp1170;
  assign tmp1170 = (tmp1167 & tmp1168) | (tmp1167 & tmp1169) | (tmp1168 & tmp1169);
  wire tmp1171;
  assign tmp1171 = (tmp1162 & tmp1166) | (tmp1162 & tmp1170) | (tmp1166 & tmp1170);
  wire tmp1172;
  assign tmp1172 = (tmp1145 & tmp1158) | (tmp1145 & tmp1171) | (tmp1158 & tmp1171);
  wire tmp1173;
  assign tmp1173 = 1'b0;
  wire tmp1174;
  assign tmp1174 = 1'b0;
  wire tmp1175;
  assign tmp1175 = 1'b0;
  wire tmp1176;
  assign tmp1176 = (tmp1173 & tmp1174) | (tmp1173 & tmp1175) | (tmp1174 & tmp1175);
  wire tmp1177;
  assign tmp1177 = 1'b0;
  wire tmp1178;
  assign tmp1178 = 1'b0;
  wire tmp1179;
  assign tmp1179 = 1'b0;
  wire tmp1180;
  assign tmp1180 = (tmp1177 & tmp1178) | (tmp1177 & tmp1179) | (tmp1178 & tmp1179);
  wire tmp1181;
  assign tmp1181 = 1'b0;
  wire tmp1182;
  assign tmp1182 = 1'b0;
  wire tmp1183;
  assign tmp1183 = 1'b0;
  wire tmp1184;
  assign tmp1184 = (tmp1181 & tmp1182) | (tmp1181 & tmp1183) | (tmp1182 & tmp1183);
  wire tmp1185;
  assign tmp1185 = (tmp1176 & tmp1180) | (tmp1176 & tmp1184) | (tmp1180 & tmp1184);
  wire tmp1186;
  assign tmp1186 = 1'b0;
  wire tmp1187;
  assign tmp1187 = 1'b0;
  wire tmp1188;
  assign tmp1188 = 1'b0;
  wire tmp1189;
  assign tmp1189 = (tmp1186 & tmp1187) | (tmp1186 & tmp1188) | (tmp1187 & tmp1188);
  wire tmp1190;
  assign tmp1190 = 1'b0;
  wire tmp1191;
  assign tmp1191 = 1'b1;
  wire tmp1192;
  assign tmp1192 = 1'b0;
  wire tmp1193;
  assign tmp1193 = (tmp1190 & tmp1191) | (tmp1190 & tmp1192) | (tmp1191 & tmp1192);
  wire tmp1194;
  assign tmp1194 = 1'b0;
  wire tmp1195;
  assign tmp1195 = 1'b0;
  wire tmp1196;
  assign tmp1196 = 1'b0;
  wire tmp1197;
  assign tmp1197 = (tmp1194 & tmp1195) | (tmp1194 & tmp1196) | (tmp1195 & tmp1196);
  wire tmp1198;
  assign tmp1198 = (tmp1189 & tmp1193) | (tmp1189 & tmp1197) | (tmp1193 & tmp1197);
  wire tmp1199;
  assign tmp1199 = 1'b0;
  wire tmp1200;
  assign tmp1200 = 1'b0;
  wire tmp1201;
  assign tmp1201 = 1'b0;
  wire tmp1202;
  assign tmp1202 = (tmp1199 & tmp1200) | (tmp1199 & tmp1201) | (tmp1200 & tmp1201);
  wire tmp1203;
  assign tmp1203 = 1'b0;
  wire tmp1204;
  assign tmp1204 = 1'b0;
  wire tmp1205;
  assign tmp1205 = 1'b0;
  wire tmp1206;
  assign tmp1206 = (tmp1203 & tmp1204) | (tmp1203 & tmp1205) | (tmp1204 & tmp1205);
  wire tmp1207;
  assign tmp1207 = 1'b0;
  wire tmp1208;
  assign tmp1208 = 1'b0;
  wire tmp1209;
  assign tmp1209 = 1'b0;
  wire tmp1210;
  assign tmp1210 = (tmp1207 & tmp1208) | (tmp1207 & tmp1209) | (tmp1208 & tmp1209);
  wire tmp1211;
  assign tmp1211 = (tmp1202 & tmp1206) | (tmp1202 & tmp1210) | (tmp1206 & tmp1210);
  wire tmp1212;
  assign tmp1212 = (tmp1185 & tmp1198) | (tmp1185 & tmp1211) | (tmp1198 & tmp1211);
  wire tmp1213;
  assign tmp1213 = (tmp1132 & tmp1172) | (tmp1132 & tmp1212) | (tmp1172 & tmp1212);
  wire tmp1214;
  assign tmp1214 = pi2;
  wire tmp1215;
  assign tmp1215 = pi3;
  wire tmp1216;
  assign tmp1216 = 1'b0;
  wire tmp1217;
  assign tmp1217 = (tmp1214 & tmp1215) | (tmp1214 & tmp1216) | (tmp1215 & tmp1216);
  wire tmp1218;
  assign tmp1218 = pi3;
  wire tmp1219;
  assign tmp1219 = 1'b1;
  wire tmp1220;
  assign tmp1220 = 1'b0;
  wire tmp1221;
  assign tmp1221 = (tmp1218 & tmp1219) | (tmp1218 & tmp1220) | (tmp1219 & tmp1220);
  wire tmp1222;
  assign tmp1222 = 1'b0;
  wire tmp1223;
  assign tmp1223 = 1'b0;
  wire tmp1224;
  assign tmp1224 = 1'b0;
  wire tmp1225;
  assign tmp1225 = (tmp1222 & tmp1223) | (tmp1222 & tmp1224) | (tmp1223 & tmp1224);
  wire tmp1226;
  assign tmp1226 = (tmp1217 & tmp1221) | (tmp1217 & tmp1225) | (tmp1221 & tmp1225);
  wire tmp1227;
  assign tmp1227 = pi3;
  wire tmp1228;
  assign tmp1228 = 1'b1;
  wire tmp1229;
  assign tmp1229 = 1'b0;
  wire tmp1230;
  assign tmp1230 = (tmp1227 & tmp1228) | (tmp1227 & tmp1229) | (tmp1228 & tmp1229);
  wire tmp1231;
  assign tmp1231 = 1'b1;
  wire tmp1232;
  assign tmp1232 = 1'b1;
  wire tmp1233;
  assign tmp1233 = 1'b1;
  wire tmp1234;
  assign tmp1234 = (tmp1231 & tmp1232) | (tmp1231 & tmp1233) | (tmp1232 & tmp1233);
  wire tmp1235;
  assign tmp1235 = 1'b0;
  wire tmp1236;
  assign tmp1236 = 1'b1;
  wire tmp1237;
  assign tmp1237 = 1'b0;
  wire tmp1238;
  assign tmp1238 = (tmp1235 & tmp1236) | (tmp1235 & tmp1237) | (tmp1236 & tmp1237);
  wire tmp1239;
  assign tmp1239 = (tmp1230 & tmp1234) | (tmp1230 & tmp1238) | (tmp1234 & tmp1238);
  wire tmp1240;
  assign tmp1240 = 1'b0;
  wire tmp1241;
  assign tmp1241 = 1'b0;
  wire tmp1242;
  assign tmp1242 = 1'b0;
  wire tmp1243;
  assign tmp1243 = (tmp1240 & tmp1241) | (tmp1240 & tmp1242) | (tmp1241 & tmp1242);
  wire tmp1244;
  assign tmp1244 = 1'b0;
  wire tmp1245;
  assign tmp1245 = 1'b1;
  wire tmp1246;
  assign tmp1246 = 1'b0;
  wire tmp1247;
  assign tmp1247 = (tmp1244 & tmp1245) | (tmp1244 & tmp1246) | (tmp1245 & tmp1246);
  wire tmp1248;
  assign tmp1248 = 1'b0;
  wire tmp1249;
  assign tmp1249 = 1'b0;
  wire tmp1250;
  assign tmp1250 = 1'b0;
  wire tmp1251;
  assign tmp1251 = (tmp1248 & tmp1249) | (tmp1248 & tmp1250) | (tmp1249 & tmp1250);
  wire tmp1252;
  assign tmp1252 = (tmp1243 & tmp1247) | (tmp1243 & tmp1251) | (tmp1247 & tmp1251);
  wire tmp1253;
  assign tmp1253 = (tmp1226 & tmp1239) | (tmp1226 & tmp1252) | (tmp1239 & tmp1252);
  wire tmp1254;
  assign tmp1254 = pi3;
  wire tmp1255;
  assign tmp1255 = 1'b1;
  wire tmp1256;
  assign tmp1256 = 1'b0;
  wire tmp1257;
  assign tmp1257 = (tmp1254 & tmp1255) | (tmp1254 & tmp1256) | (tmp1255 & tmp1256);
  wire tmp1258;
  assign tmp1258 = 1'b1;
  wire tmp1259;
  assign tmp1259 = 1'b1;
  wire tmp1260;
  assign tmp1260 = 1'b1;
  wire tmp1261;
  assign tmp1261 = (tmp1258 & tmp1259) | (tmp1258 & tmp1260) | (tmp1259 & tmp1260);
  wire tmp1262;
  assign tmp1262 = 1'b0;
  wire tmp1263;
  assign tmp1263 = 1'b1;
  wire tmp1264;
  assign tmp1264 = 1'b0;
  wire tmp1265;
  assign tmp1265 = (tmp1262 & tmp1263) | (tmp1262 & tmp1264) | (tmp1263 & tmp1264);
  wire tmp1266;
  assign tmp1266 = (tmp1257 & tmp1261) | (tmp1257 & tmp1265) | (tmp1261 & tmp1265);
  wire tmp1267;
  assign tmp1267 = 1'b1;
  wire tmp1268;
  assign tmp1268 = 1'b1;
  wire tmp1269;
  assign tmp1269 = 1'b1;
  wire tmp1270;
  assign tmp1270 = (tmp1267 & tmp1268) | (tmp1267 & tmp1269) | (tmp1268 & tmp1269);
  wire tmp1271;
  assign tmp1271 = 1'b1;
  wire tmp1272;
  assign tmp1272 = 1'b1;
  wire tmp1273;
  assign tmp1273 = 1'b1;
  wire tmp1274;
  assign tmp1274 = (tmp1271 & tmp1272) | (tmp1271 & tmp1273) | (tmp1272 & tmp1273);
  wire tmp1275;
  assign tmp1275 = 1'b1;
  wire tmp1276;
  assign tmp1276 = 1'b1;
  wire tmp1277;
  assign tmp1277 = 1'b1;
  wire tmp1278;
  assign tmp1278 = (tmp1275 & tmp1276) | (tmp1275 & tmp1277) | (tmp1276 & tmp1277);
  wire tmp1279;
  assign tmp1279 = (tmp1270 & tmp1274) | (tmp1270 & tmp1278) | (tmp1274 & tmp1278);
  wire tmp1280;
  assign tmp1280 = 1'b0;
  wire tmp1281;
  assign tmp1281 = 1'b1;
  wire tmp1282;
  assign tmp1282 = 1'b0;
  wire tmp1283;
  assign tmp1283 = (tmp1280 & tmp1281) | (tmp1280 & tmp1282) | (tmp1281 & tmp1282);
  wire tmp1284;
  assign tmp1284 = 1'b1;
  wire tmp1285;
  assign tmp1285 = 1'b1;
  wire tmp1286;
  assign tmp1286 = 1'b1;
  wire tmp1287;
  assign tmp1287 = (tmp1284 & tmp1285) | (tmp1284 & tmp1286) | (tmp1285 & tmp1286);
  wire tmp1288;
  assign tmp1288 = 1'b0;
  wire tmp1289;
  assign tmp1289 = 1'b1;
  wire tmp1290;
  assign tmp1290 = 1'b0;
  wire tmp1291;
  assign tmp1291 = (tmp1288 & tmp1289) | (tmp1288 & tmp1290) | (tmp1289 & tmp1290);
  wire tmp1292;
  assign tmp1292 = (tmp1283 & tmp1287) | (tmp1283 & tmp1291) | (tmp1287 & tmp1291);
  wire tmp1293;
  assign tmp1293 = (tmp1266 & tmp1279) | (tmp1266 & tmp1292) | (tmp1279 & tmp1292);
  wire tmp1294;
  assign tmp1294 = 1'b0;
  wire tmp1295;
  assign tmp1295 = 1'b0;
  wire tmp1296;
  assign tmp1296 = 1'b0;
  wire tmp1297;
  assign tmp1297 = (tmp1294 & tmp1295) | (tmp1294 & tmp1296) | (tmp1295 & tmp1296);
  wire tmp1298;
  assign tmp1298 = 1'b0;
  wire tmp1299;
  assign tmp1299 = 1'b1;
  wire tmp1300;
  assign tmp1300 = 1'b0;
  wire tmp1301;
  assign tmp1301 = (tmp1298 & tmp1299) | (tmp1298 & tmp1300) | (tmp1299 & tmp1300);
  wire tmp1302;
  assign tmp1302 = 1'b0;
  wire tmp1303;
  assign tmp1303 = 1'b0;
  wire tmp1304;
  assign tmp1304 = 1'b0;
  wire tmp1305;
  assign tmp1305 = (tmp1302 & tmp1303) | (tmp1302 & tmp1304) | (tmp1303 & tmp1304);
  wire tmp1306;
  assign tmp1306 = (tmp1297 & tmp1301) | (tmp1297 & tmp1305) | (tmp1301 & tmp1305);
  wire tmp1307;
  assign tmp1307 = 1'b0;
  wire tmp1308;
  assign tmp1308 = 1'b1;
  wire tmp1309;
  assign tmp1309 = 1'b0;
  wire tmp1310;
  assign tmp1310 = (tmp1307 & tmp1308) | (tmp1307 & tmp1309) | (tmp1308 & tmp1309);
  wire tmp1311;
  assign tmp1311 = 1'b1;
  wire tmp1312;
  assign tmp1312 = 1'b1;
  wire tmp1313;
  assign tmp1313 = 1'b1;
  wire tmp1314;
  assign tmp1314 = (tmp1311 & tmp1312) | (tmp1311 & tmp1313) | (tmp1312 & tmp1313);
  wire tmp1315;
  assign tmp1315 = 1'b0;
  wire tmp1316;
  assign tmp1316 = 1'b1;
  wire tmp1317;
  assign tmp1317 = 1'b0;
  wire tmp1318;
  assign tmp1318 = (tmp1315 & tmp1316) | (tmp1315 & tmp1317) | (tmp1316 & tmp1317);
  wire tmp1319;
  assign tmp1319 = (tmp1310 & tmp1314) | (tmp1310 & tmp1318) | (tmp1314 & tmp1318);
  wire tmp1320;
  assign tmp1320 = 1'b0;
  wire tmp1321;
  assign tmp1321 = 1'b0;
  wire tmp1322;
  assign tmp1322 = 1'b0;
  wire tmp1323;
  assign tmp1323 = (tmp1320 & tmp1321) | (tmp1320 & tmp1322) | (tmp1321 & tmp1322);
  wire tmp1324;
  assign tmp1324 = 1'b0;
  wire tmp1325;
  assign tmp1325 = 1'b1;
  wire tmp1326;
  assign tmp1326 = 1'b0;
  wire tmp1327;
  assign tmp1327 = (tmp1324 & tmp1325) | (tmp1324 & tmp1326) | (tmp1325 & tmp1326);
  wire tmp1328;
  assign tmp1328 = 1'b0;
  wire tmp1329;
  assign tmp1329 = 1'b0;
  wire tmp1330;
  assign tmp1330 = 1'b0;
  wire tmp1331;
  assign tmp1331 = (tmp1328 & tmp1329) | (tmp1328 & tmp1330) | (tmp1329 & tmp1330);
  wire tmp1332;
  assign tmp1332 = (tmp1323 & tmp1327) | (tmp1323 & tmp1331) | (tmp1327 & tmp1331);
  wire tmp1333;
  assign tmp1333 = (tmp1306 & tmp1319) | (tmp1306 & tmp1332) | (tmp1319 & tmp1332);
  wire tmp1334;
  assign tmp1334 = (tmp1253 & tmp1293) | (tmp1253 & tmp1333) | (tmp1293 & tmp1333);
  wire tmp1335;
  assign tmp1335 = 1'b0;
  wire tmp1336;
  assign tmp1336 = 1'b0;
  wire tmp1337;
  assign tmp1337 = 1'b0;
  wire tmp1338;
  assign tmp1338 = (tmp1335 & tmp1336) | (tmp1335 & tmp1337) | (tmp1336 & tmp1337);
  wire tmp1339;
  assign tmp1339 = 1'b0;
  wire tmp1340;
  assign tmp1340 = 1'b0;
  wire tmp1341;
  assign tmp1341 = 1'b0;
  wire tmp1342;
  assign tmp1342 = (tmp1339 & tmp1340) | (tmp1339 & tmp1341) | (tmp1340 & tmp1341);
  wire tmp1343;
  assign tmp1343 = 1'b0;
  wire tmp1344;
  assign tmp1344 = 1'b0;
  wire tmp1345;
  assign tmp1345 = 1'b0;
  wire tmp1346;
  assign tmp1346 = (tmp1343 & tmp1344) | (tmp1343 & tmp1345) | (tmp1344 & tmp1345);
  wire tmp1347;
  assign tmp1347 = (tmp1338 & tmp1342) | (tmp1338 & tmp1346) | (tmp1342 & tmp1346);
  wire tmp1348;
  assign tmp1348 = 1'b0;
  wire tmp1349;
  assign tmp1349 = 1'b0;
  wire tmp1350;
  assign tmp1350 = 1'b0;
  wire tmp1351;
  assign tmp1351 = (tmp1348 & tmp1349) | (tmp1348 & tmp1350) | (tmp1349 & tmp1350);
  wire tmp1352;
  assign tmp1352 = 1'b0;
  wire tmp1353;
  assign tmp1353 = 1'b1;
  wire tmp1354;
  assign tmp1354 = 1'b0;
  wire tmp1355;
  assign tmp1355 = (tmp1352 & tmp1353) | (tmp1352 & tmp1354) | (tmp1353 & tmp1354);
  wire tmp1356;
  assign tmp1356 = 1'b0;
  wire tmp1357;
  assign tmp1357 = 1'b0;
  wire tmp1358;
  assign tmp1358 = 1'b0;
  wire tmp1359;
  assign tmp1359 = (tmp1356 & tmp1357) | (tmp1356 & tmp1358) | (tmp1357 & tmp1358);
  wire tmp1360;
  assign tmp1360 = (tmp1351 & tmp1355) | (tmp1351 & tmp1359) | (tmp1355 & tmp1359);
  wire tmp1361;
  assign tmp1361 = 1'b0;
  wire tmp1362;
  assign tmp1362 = 1'b0;
  wire tmp1363;
  assign tmp1363 = 1'b0;
  wire tmp1364;
  assign tmp1364 = (tmp1361 & tmp1362) | (tmp1361 & tmp1363) | (tmp1362 & tmp1363);
  wire tmp1365;
  assign tmp1365 = 1'b0;
  wire tmp1366;
  assign tmp1366 = 1'b0;
  wire tmp1367;
  assign tmp1367 = 1'b0;
  wire tmp1368;
  assign tmp1368 = (tmp1365 & tmp1366) | (tmp1365 & tmp1367) | (tmp1366 & tmp1367);
  wire tmp1369;
  assign tmp1369 = 1'b0;
  wire tmp1370;
  assign tmp1370 = 1'b0;
  wire tmp1371;
  assign tmp1371 = 1'b0;
  wire tmp1372;
  assign tmp1372 = (tmp1369 & tmp1370) | (tmp1369 & tmp1371) | (tmp1370 & tmp1371);
  wire tmp1373;
  assign tmp1373 = (tmp1364 & tmp1368) | (tmp1364 & tmp1372) | (tmp1368 & tmp1372);
  wire tmp1374;
  assign tmp1374 = (tmp1347 & tmp1360) | (tmp1347 & tmp1373) | (tmp1360 & tmp1373);
  wire tmp1375;
  assign tmp1375 = 1'b0;
  wire tmp1376;
  assign tmp1376 = 1'b0;
  wire tmp1377;
  assign tmp1377 = 1'b0;
  wire tmp1378;
  assign tmp1378 = (tmp1375 & tmp1376) | (tmp1375 & tmp1377) | (tmp1376 & tmp1377);
  wire tmp1379;
  assign tmp1379 = 1'b0;
  wire tmp1380;
  assign tmp1380 = 1'b1;
  wire tmp1381;
  assign tmp1381 = 1'b0;
  wire tmp1382;
  assign tmp1382 = (tmp1379 & tmp1380) | (tmp1379 & tmp1381) | (tmp1380 & tmp1381);
  wire tmp1383;
  assign tmp1383 = 1'b0;
  wire tmp1384;
  assign tmp1384 = 1'b0;
  wire tmp1385;
  assign tmp1385 = 1'b0;
  wire tmp1386;
  assign tmp1386 = (tmp1383 & tmp1384) | (tmp1383 & tmp1385) | (tmp1384 & tmp1385);
  wire tmp1387;
  assign tmp1387 = (tmp1378 & tmp1382) | (tmp1378 & tmp1386) | (tmp1382 & tmp1386);
  wire tmp1388;
  assign tmp1388 = 1'b0;
  wire tmp1389;
  assign tmp1389 = 1'b1;
  wire tmp1390;
  assign tmp1390 = 1'b0;
  wire tmp1391;
  assign tmp1391 = (tmp1388 & tmp1389) | (tmp1388 & tmp1390) | (tmp1389 & tmp1390);
  wire tmp1392;
  assign tmp1392 = 1'b1;
  wire tmp1393;
  assign tmp1393 = 1'b1;
  wire tmp1394;
  assign tmp1394 = 1'b1;
  wire tmp1395;
  assign tmp1395 = (tmp1392 & tmp1393) | (tmp1392 & tmp1394) | (tmp1393 & tmp1394);
  wire tmp1396;
  assign tmp1396 = 1'b0;
  wire tmp1397;
  assign tmp1397 = 1'b1;
  wire tmp1398;
  assign tmp1398 = 1'b0;
  wire tmp1399;
  assign tmp1399 = (tmp1396 & tmp1397) | (tmp1396 & tmp1398) | (tmp1397 & tmp1398);
  wire tmp1400;
  assign tmp1400 = (tmp1391 & tmp1395) | (tmp1391 & tmp1399) | (tmp1395 & tmp1399);
  wire tmp1401;
  assign tmp1401 = 1'b0;
  wire tmp1402;
  assign tmp1402 = 1'b0;
  wire tmp1403;
  assign tmp1403 = 1'b0;
  wire tmp1404;
  assign tmp1404 = (tmp1401 & tmp1402) | (tmp1401 & tmp1403) | (tmp1402 & tmp1403);
  wire tmp1405;
  assign tmp1405 = 1'b0;
  wire tmp1406;
  assign tmp1406 = 1'b1;
  wire tmp1407;
  assign tmp1407 = 1'b0;
  wire tmp1408;
  assign tmp1408 = (tmp1405 & tmp1406) | (tmp1405 & tmp1407) | (tmp1406 & tmp1407);
  wire tmp1409;
  assign tmp1409 = 1'b0;
  wire tmp1410;
  assign tmp1410 = 1'b0;
  wire tmp1411;
  assign tmp1411 = 1'b0;
  wire tmp1412;
  assign tmp1412 = (tmp1409 & tmp1410) | (tmp1409 & tmp1411) | (tmp1410 & tmp1411);
  wire tmp1413;
  assign tmp1413 = (tmp1404 & tmp1408) | (tmp1404 & tmp1412) | (tmp1408 & tmp1412);
  wire tmp1414;
  assign tmp1414 = (tmp1387 & tmp1400) | (tmp1387 & tmp1413) | (tmp1400 & tmp1413);
  wire tmp1415;
  assign tmp1415 = 1'b0;
  wire tmp1416;
  assign tmp1416 = 1'b0;
  wire tmp1417;
  assign tmp1417 = 1'b0;
  wire tmp1418;
  assign tmp1418 = (tmp1415 & tmp1416) | (tmp1415 & tmp1417) | (tmp1416 & tmp1417);
  wire tmp1419;
  assign tmp1419 = 1'b0;
  wire tmp1420;
  assign tmp1420 = 1'b0;
  wire tmp1421;
  assign tmp1421 = 1'b0;
  wire tmp1422;
  assign tmp1422 = (tmp1419 & tmp1420) | (tmp1419 & tmp1421) | (tmp1420 & tmp1421);
  wire tmp1423;
  assign tmp1423 = 1'b0;
  wire tmp1424;
  assign tmp1424 = 1'b0;
  wire tmp1425;
  assign tmp1425 = 1'b0;
  wire tmp1426;
  assign tmp1426 = (tmp1423 & tmp1424) | (tmp1423 & tmp1425) | (tmp1424 & tmp1425);
  wire tmp1427;
  assign tmp1427 = (tmp1418 & tmp1422) | (tmp1418 & tmp1426) | (tmp1422 & tmp1426);
  wire tmp1428;
  assign tmp1428 = 1'b0;
  wire tmp1429;
  assign tmp1429 = 1'b0;
  wire tmp1430;
  assign tmp1430 = 1'b0;
  wire tmp1431;
  assign tmp1431 = (tmp1428 & tmp1429) | (tmp1428 & tmp1430) | (tmp1429 & tmp1430);
  wire tmp1432;
  assign tmp1432 = 1'b0;
  wire tmp1433;
  assign tmp1433 = 1'b1;
  wire tmp1434;
  assign tmp1434 = 1'b0;
  wire tmp1435;
  assign tmp1435 = (tmp1432 & tmp1433) | (tmp1432 & tmp1434) | (tmp1433 & tmp1434);
  wire tmp1436;
  assign tmp1436 = 1'b0;
  wire tmp1437;
  assign tmp1437 = 1'b0;
  wire tmp1438;
  assign tmp1438 = 1'b0;
  wire tmp1439;
  assign tmp1439 = (tmp1436 & tmp1437) | (tmp1436 & tmp1438) | (tmp1437 & tmp1438);
  wire tmp1440;
  assign tmp1440 = (tmp1431 & tmp1435) | (tmp1431 & tmp1439) | (tmp1435 & tmp1439);
  wire tmp1441;
  assign tmp1441 = 1'b0;
  wire tmp1442;
  assign tmp1442 = 1'b0;
  wire tmp1443;
  assign tmp1443 = 1'b0;
  wire tmp1444;
  assign tmp1444 = (tmp1441 & tmp1442) | (tmp1441 & tmp1443) | (tmp1442 & tmp1443);
  wire tmp1445;
  assign tmp1445 = 1'b0;
  wire tmp1446;
  assign tmp1446 = 1'b0;
  wire tmp1447;
  assign tmp1447 = 1'b0;
  wire tmp1448;
  assign tmp1448 = (tmp1445 & tmp1446) | (tmp1445 & tmp1447) | (tmp1446 & tmp1447);
  wire tmp1449;
  assign tmp1449 = 1'b0;
  wire tmp1450;
  assign tmp1450 = 1'b0;
  wire tmp1451;
  assign tmp1451 = 1'b0;
  wire tmp1452;
  assign tmp1452 = (tmp1449 & tmp1450) | (tmp1449 & tmp1451) | (tmp1450 & tmp1451);
  wire tmp1453;
  assign tmp1453 = (tmp1444 & tmp1448) | (tmp1444 & tmp1452) | (tmp1448 & tmp1452);
  wire tmp1454;
  assign tmp1454 = (tmp1427 & tmp1440) | (tmp1427 & tmp1453) | (tmp1440 & tmp1453);
  wire tmp1455;
  assign tmp1455 = (tmp1374 & tmp1414) | (tmp1374 & tmp1454) | (tmp1414 & tmp1454);
  wire tmp1456;
  assign tmp1456 = (tmp1213 & tmp1334) | (tmp1213 & tmp1455) | (tmp1334 & tmp1455);
  wire tmp1457;
  assign tmp1457 = pi2;
  wire tmp1458;
  assign tmp1458 = pi3;
  wire tmp1459;
  assign tmp1459 = 1'b0;
  wire tmp1460;
  assign tmp1460 = (tmp1457 & tmp1458) | (tmp1457 & tmp1459) | (tmp1458 & tmp1459);
  wire tmp1461;
  assign tmp1461 = pi3;
  wire tmp1462;
  assign tmp1462 = 1'b1;
  wire tmp1463;
  assign tmp1463 = 1'b0;
  wire tmp1464;
  assign tmp1464 = (tmp1461 & tmp1462) | (tmp1461 & tmp1463) | (tmp1462 & tmp1463);
  wire tmp1465;
  assign tmp1465 = 1'b0;
  wire tmp1466;
  assign tmp1466 = 1'b0;
  wire tmp1467;
  assign tmp1467 = 1'b0;
  wire tmp1468;
  assign tmp1468 = (tmp1465 & tmp1466) | (tmp1465 & tmp1467) | (tmp1466 & tmp1467);
  wire tmp1469;
  assign tmp1469 = (tmp1460 & tmp1464) | (tmp1460 & tmp1468) | (tmp1464 & tmp1468);
  wire tmp1470;
  assign tmp1470 = pi3;
  wire tmp1471;
  assign tmp1471 = 1'b1;
  wire tmp1472;
  assign tmp1472 = 1'b0;
  wire tmp1473;
  assign tmp1473 = (tmp1470 & tmp1471) | (tmp1470 & tmp1472) | (tmp1471 & tmp1472);
  wire tmp1474;
  assign tmp1474 = 1'b1;
  wire tmp1475;
  assign tmp1475 = 1'b1;
  wire tmp1476;
  assign tmp1476 = 1'b1;
  wire tmp1477;
  assign tmp1477 = (tmp1474 & tmp1475) | (tmp1474 & tmp1476) | (tmp1475 & tmp1476);
  wire tmp1478;
  assign tmp1478 = 1'b0;
  wire tmp1479;
  assign tmp1479 = 1'b1;
  wire tmp1480;
  assign tmp1480 = 1'b0;
  wire tmp1481;
  assign tmp1481 = (tmp1478 & tmp1479) | (tmp1478 & tmp1480) | (tmp1479 & tmp1480);
  wire tmp1482;
  assign tmp1482 = (tmp1473 & tmp1477) | (tmp1473 & tmp1481) | (tmp1477 & tmp1481);
  wire tmp1483;
  assign tmp1483 = 1'b0;
  wire tmp1484;
  assign tmp1484 = 1'b0;
  wire tmp1485;
  assign tmp1485 = 1'b0;
  wire tmp1486;
  assign tmp1486 = (tmp1483 & tmp1484) | (tmp1483 & tmp1485) | (tmp1484 & tmp1485);
  wire tmp1487;
  assign tmp1487 = 1'b0;
  wire tmp1488;
  assign tmp1488 = 1'b1;
  wire tmp1489;
  assign tmp1489 = 1'b0;
  wire tmp1490;
  assign tmp1490 = (tmp1487 & tmp1488) | (tmp1487 & tmp1489) | (tmp1488 & tmp1489);
  wire tmp1491;
  assign tmp1491 = 1'b0;
  wire tmp1492;
  assign tmp1492 = 1'b0;
  wire tmp1493;
  assign tmp1493 = 1'b0;
  wire tmp1494;
  assign tmp1494 = (tmp1491 & tmp1492) | (tmp1491 & tmp1493) | (tmp1492 & tmp1493);
  wire tmp1495;
  assign tmp1495 = (tmp1486 & tmp1490) | (tmp1486 & tmp1494) | (tmp1490 & tmp1494);
  wire tmp1496;
  assign tmp1496 = (tmp1469 & tmp1482) | (tmp1469 & tmp1495) | (tmp1482 & tmp1495);
  wire tmp1497;
  assign tmp1497 = pi3;
  wire tmp1498;
  assign tmp1498 = 1'b1;
  wire tmp1499;
  assign tmp1499 = 1'b0;
  wire tmp1500;
  assign tmp1500 = (tmp1497 & tmp1498) | (tmp1497 & tmp1499) | (tmp1498 & tmp1499);
  wire tmp1501;
  assign tmp1501 = 1'b1;
  wire tmp1502;
  assign tmp1502 = 1'b1;
  wire tmp1503;
  assign tmp1503 = 1'b1;
  wire tmp1504;
  assign tmp1504 = (tmp1501 & tmp1502) | (tmp1501 & tmp1503) | (tmp1502 & tmp1503);
  wire tmp1505;
  assign tmp1505 = 1'b0;
  wire tmp1506;
  assign tmp1506 = 1'b1;
  wire tmp1507;
  assign tmp1507 = 1'b0;
  wire tmp1508;
  assign tmp1508 = (tmp1505 & tmp1506) | (tmp1505 & tmp1507) | (tmp1506 & tmp1507);
  wire tmp1509;
  assign tmp1509 = (tmp1500 & tmp1504) | (tmp1500 & tmp1508) | (tmp1504 & tmp1508);
  wire tmp1510;
  assign tmp1510 = 1'b1;
  wire tmp1511;
  assign tmp1511 = 1'b1;
  wire tmp1512;
  assign tmp1512 = 1'b1;
  wire tmp1513;
  assign tmp1513 = (tmp1510 & tmp1511) | (tmp1510 & tmp1512) | (tmp1511 & tmp1512);
  wire tmp1514;
  assign tmp1514 = 1'b1;
  wire tmp1515;
  assign tmp1515 = 1'b1;
  wire tmp1516;
  assign tmp1516 = 1'b1;
  wire tmp1517;
  assign tmp1517 = (tmp1514 & tmp1515) | (tmp1514 & tmp1516) | (tmp1515 & tmp1516);
  wire tmp1518;
  assign tmp1518 = 1'b1;
  wire tmp1519;
  assign tmp1519 = 1'b1;
  wire tmp1520;
  assign tmp1520 = 1'b1;
  wire tmp1521;
  assign tmp1521 = (tmp1518 & tmp1519) | (tmp1518 & tmp1520) | (tmp1519 & tmp1520);
  wire tmp1522;
  assign tmp1522 = (tmp1513 & tmp1517) | (tmp1513 & tmp1521) | (tmp1517 & tmp1521);
  wire tmp1523;
  assign tmp1523 = 1'b0;
  wire tmp1524;
  assign tmp1524 = 1'b1;
  wire tmp1525;
  assign tmp1525 = 1'b0;
  wire tmp1526;
  assign tmp1526 = (tmp1523 & tmp1524) | (tmp1523 & tmp1525) | (tmp1524 & tmp1525);
  wire tmp1527;
  assign tmp1527 = 1'b1;
  wire tmp1528;
  assign tmp1528 = 1'b1;
  wire tmp1529;
  assign tmp1529 = 1'b1;
  wire tmp1530;
  assign tmp1530 = (tmp1527 & tmp1528) | (tmp1527 & tmp1529) | (tmp1528 & tmp1529);
  wire tmp1531;
  assign tmp1531 = 1'b0;
  wire tmp1532;
  assign tmp1532 = 1'b1;
  wire tmp1533;
  assign tmp1533 = 1'b0;
  wire tmp1534;
  assign tmp1534 = (tmp1531 & tmp1532) | (tmp1531 & tmp1533) | (tmp1532 & tmp1533);
  wire tmp1535;
  assign tmp1535 = (tmp1526 & tmp1530) | (tmp1526 & tmp1534) | (tmp1530 & tmp1534);
  wire tmp1536;
  assign tmp1536 = (tmp1509 & tmp1522) | (tmp1509 & tmp1535) | (tmp1522 & tmp1535);
  wire tmp1537;
  assign tmp1537 = 1'b0;
  wire tmp1538;
  assign tmp1538 = 1'b0;
  wire tmp1539;
  assign tmp1539 = 1'b0;
  wire tmp1540;
  assign tmp1540 = (tmp1537 & tmp1538) | (tmp1537 & tmp1539) | (tmp1538 & tmp1539);
  wire tmp1541;
  assign tmp1541 = 1'b0;
  wire tmp1542;
  assign tmp1542 = 1'b1;
  wire tmp1543;
  assign tmp1543 = 1'b0;
  wire tmp1544;
  assign tmp1544 = (tmp1541 & tmp1542) | (tmp1541 & tmp1543) | (tmp1542 & tmp1543);
  wire tmp1545;
  assign tmp1545 = 1'b0;
  wire tmp1546;
  assign tmp1546 = 1'b0;
  wire tmp1547;
  assign tmp1547 = 1'b0;
  wire tmp1548;
  assign tmp1548 = (tmp1545 & tmp1546) | (tmp1545 & tmp1547) | (tmp1546 & tmp1547);
  wire tmp1549;
  assign tmp1549 = (tmp1540 & tmp1544) | (tmp1540 & tmp1548) | (tmp1544 & tmp1548);
  wire tmp1550;
  assign tmp1550 = 1'b0;
  wire tmp1551;
  assign tmp1551 = 1'b1;
  wire tmp1552;
  assign tmp1552 = 1'b0;
  wire tmp1553;
  assign tmp1553 = (tmp1550 & tmp1551) | (tmp1550 & tmp1552) | (tmp1551 & tmp1552);
  wire tmp1554;
  assign tmp1554 = 1'b1;
  wire tmp1555;
  assign tmp1555 = 1'b1;
  wire tmp1556;
  assign tmp1556 = 1'b1;
  wire tmp1557;
  assign tmp1557 = (tmp1554 & tmp1555) | (tmp1554 & tmp1556) | (tmp1555 & tmp1556);
  wire tmp1558;
  assign tmp1558 = 1'b0;
  wire tmp1559;
  assign tmp1559 = 1'b1;
  wire tmp1560;
  assign tmp1560 = 1'b0;
  wire tmp1561;
  assign tmp1561 = (tmp1558 & tmp1559) | (tmp1558 & tmp1560) | (tmp1559 & tmp1560);
  wire tmp1562;
  assign tmp1562 = (tmp1553 & tmp1557) | (tmp1553 & tmp1561) | (tmp1557 & tmp1561);
  wire tmp1563;
  assign tmp1563 = 1'b0;
  wire tmp1564;
  assign tmp1564 = 1'b0;
  wire tmp1565;
  assign tmp1565 = 1'b0;
  wire tmp1566;
  assign tmp1566 = (tmp1563 & tmp1564) | (tmp1563 & tmp1565) | (tmp1564 & tmp1565);
  wire tmp1567;
  assign tmp1567 = 1'b0;
  wire tmp1568;
  assign tmp1568 = 1'b1;
  wire tmp1569;
  assign tmp1569 = 1'b0;
  wire tmp1570;
  assign tmp1570 = (tmp1567 & tmp1568) | (tmp1567 & tmp1569) | (tmp1568 & tmp1569);
  wire tmp1571;
  assign tmp1571 = 1'b0;
  wire tmp1572;
  assign tmp1572 = 1'b0;
  wire tmp1573;
  assign tmp1573 = 1'b0;
  wire tmp1574;
  assign tmp1574 = (tmp1571 & tmp1572) | (tmp1571 & tmp1573) | (tmp1572 & tmp1573);
  wire tmp1575;
  assign tmp1575 = (tmp1566 & tmp1570) | (tmp1566 & tmp1574) | (tmp1570 & tmp1574);
  wire tmp1576;
  assign tmp1576 = (tmp1549 & tmp1562) | (tmp1549 & tmp1575) | (tmp1562 & tmp1575);
  wire tmp1577;
  assign tmp1577 = (tmp1496 & tmp1536) | (tmp1496 & tmp1576) | (tmp1536 & tmp1576);
  wire tmp1578;
  assign tmp1578 = pi3;
  wire tmp1579;
  assign tmp1579 = 1'b1;
  wire tmp1580;
  assign tmp1580 = 1'b0;
  wire tmp1581;
  assign tmp1581 = (tmp1578 & tmp1579) | (tmp1578 & tmp1580) | (tmp1579 & tmp1580);
  wire tmp1582;
  assign tmp1582 = 1'b1;
  wire tmp1583;
  assign tmp1583 = 1'b1;
  wire tmp1584;
  assign tmp1584 = 1'b1;
  wire tmp1585;
  assign tmp1585 = (tmp1582 & tmp1583) | (tmp1582 & tmp1584) | (tmp1583 & tmp1584);
  wire tmp1586;
  assign tmp1586 = 1'b0;
  wire tmp1587;
  assign tmp1587 = 1'b1;
  wire tmp1588;
  assign tmp1588 = 1'b0;
  wire tmp1589;
  assign tmp1589 = (tmp1586 & tmp1587) | (tmp1586 & tmp1588) | (tmp1587 & tmp1588);
  wire tmp1590;
  assign tmp1590 = (tmp1581 & tmp1585) | (tmp1581 & tmp1589) | (tmp1585 & tmp1589);
  wire tmp1591;
  assign tmp1591 = 1'b1;
  wire tmp1592;
  assign tmp1592 = 1'b1;
  wire tmp1593;
  assign tmp1593 = 1'b1;
  wire tmp1594;
  assign tmp1594 = (tmp1591 & tmp1592) | (tmp1591 & tmp1593) | (tmp1592 & tmp1593);
  wire tmp1595;
  assign tmp1595 = 1'b1;
  wire tmp1596;
  assign tmp1596 = 1'b1;
  wire tmp1597;
  assign tmp1597 = 1'b1;
  wire tmp1598;
  assign tmp1598 = (tmp1595 & tmp1596) | (tmp1595 & tmp1597) | (tmp1596 & tmp1597);
  wire tmp1599;
  assign tmp1599 = 1'b1;
  wire tmp1600;
  assign tmp1600 = 1'b1;
  wire tmp1601;
  assign tmp1601 = 1'b1;
  wire tmp1602;
  assign tmp1602 = (tmp1599 & tmp1600) | (tmp1599 & tmp1601) | (tmp1600 & tmp1601);
  wire tmp1603;
  assign tmp1603 = (tmp1594 & tmp1598) | (tmp1594 & tmp1602) | (tmp1598 & tmp1602);
  wire tmp1604;
  assign tmp1604 = 1'b0;
  wire tmp1605;
  assign tmp1605 = 1'b1;
  wire tmp1606;
  assign tmp1606 = 1'b0;
  wire tmp1607;
  assign tmp1607 = (tmp1604 & tmp1605) | (tmp1604 & tmp1606) | (tmp1605 & tmp1606);
  wire tmp1608;
  assign tmp1608 = 1'b1;
  wire tmp1609;
  assign tmp1609 = 1'b1;
  wire tmp1610;
  assign tmp1610 = 1'b1;
  wire tmp1611;
  assign tmp1611 = (tmp1608 & tmp1609) | (tmp1608 & tmp1610) | (tmp1609 & tmp1610);
  wire tmp1612;
  assign tmp1612 = 1'b0;
  wire tmp1613;
  assign tmp1613 = 1'b1;
  wire tmp1614;
  assign tmp1614 = 1'b0;
  wire tmp1615;
  assign tmp1615 = (tmp1612 & tmp1613) | (tmp1612 & tmp1614) | (tmp1613 & tmp1614);
  wire tmp1616;
  assign tmp1616 = (tmp1607 & tmp1611) | (tmp1607 & tmp1615) | (tmp1611 & tmp1615);
  wire tmp1617;
  assign tmp1617 = (tmp1590 & tmp1603) | (tmp1590 & tmp1616) | (tmp1603 & tmp1616);
  wire tmp1618;
  assign tmp1618 = 1'b1;
  wire tmp1619;
  assign tmp1619 = 1'b1;
  wire tmp1620;
  assign tmp1620 = 1'b1;
  wire tmp1621;
  assign tmp1621 = (tmp1618 & tmp1619) | (tmp1618 & tmp1620) | (tmp1619 & tmp1620);
  wire tmp1622;
  assign tmp1622 = 1'b1;
  wire tmp1623;
  assign tmp1623 = 1'b1;
  wire tmp1624;
  assign tmp1624 = 1'b1;
  wire tmp1625;
  assign tmp1625 = (tmp1622 & tmp1623) | (tmp1622 & tmp1624) | (tmp1623 & tmp1624);
  wire tmp1626;
  assign tmp1626 = 1'b1;
  wire tmp1627;
  assign tmp1627 = 1'b1;
  wire tmp1628;
  assign tmp1628 = 1'b1;
  wire tmp1629;
  assign tmp1629 = (tmp1626 & tmp1627) | (tmp1626 & tmp1628) | (tmp1627 & tmp1628);
  wire tmp1630;
  assign tmp1630 = (tmp1621 & tmp1625) | (tmp1621 & tmp1629) | (tmp1625 & tmp1629);
  wire tmp1631;
  assign tmp1631 = 1'b1;
  wire tmp1632;
  assign tmp1632 = 1'b1;
  wire tmp1633;
  assign tmp1633 = 1'b1;
  wire tmp1634;
  assign tmp1634 = (tmp1631 & tmp1632) | (tmp1631 & tmp1633) | (tmp1632 & tmp1633);
  wire tmp1635;
  assign tmp1635 = 1'b1;
  wire tmp1636;
  assign tmp1636 = ~pi4;
  wire tmp1637;
  assign tmp1637 = ~pi5;
  wire tmp1638;
  assign tmp1638 = (tmp1635 & tmp1636) | (tmp1635 & tmp1637) | (tmp1636 & tmp1637);
  wire tmp1639;
  assign tmp1639 = 1'b1;
  wire tmp1640;
  assign tmp1640 = ~pi5;
  wire tmp1641;
  assign tmp1641 = ~pi6;
  wire tmp1642;
  assign tmp1642 = (tmp1639 & tmp1640) | (tmp1639 & tmp1641) | (tmp1640 & tmp1641);
  wire tmp1643;
  assign tmp1643 = (tmp1634 & tmp1638) | (tmp1634 & tmp1642) | (tmp1638 & tmp1642);
  wire tmp1644;
  assign tmp1644 = 1'b1;
  wire tmp1645;
  assign tmp1645 = 1'b1;
  wire tmp1646;
  assign tmp1646 = 1'b1;
  wire tmp1647;
  assign tmp1647 = (tmp1644 & tmp1645) | (tmp1644 & tmp1646) | (tmp1645 & tmp1646);
  wire tmp1648;
  assign tmp1648 = 1'b1;
  wire tmp1649;
  assign tmp1649 = ~pi5;
  wire tmp1650;
  assign tmp1650 = ~pi6;
  wire tmp1651;
  assign tmp1651 = (tmp1648 & tmp1649) | (tmp1648 & tmp1650) | (tmp1649 & tmp1650);
  wire tmp1652;
  assign tmp1652 = 1'b1;
  wire tmp1653;
  assign tmp1653 = ~pi6;
  wire tmp1654;
  assign tmp1654 = ~pi7;
  wire tmp1655;
  assign tmp1655 = (tmp1652 & tmp1653) | (tmp1652 & tmp1654) | (tmp1653 & tmp1654);
  wire tmp1656;
  assign tmp1656 = (tmp1647 & tmp1651) | (tmp1647 & tmp1655) | (tmp1651 & tmp1655);
  wire tmp1657;
  assign tmp1657 = (tmp1630 & tmp1643) | (tmp1630 & tmp1656) | (tmp1643 & tmp1656);
  wire tmp1658;
  assign tmp1658 = 1'b0;
  wire tmp1659;
  assign tmp1659 = 1'b1;
  wire tmp1660;
  assign tmp1660 = 1'b0;
  wire tmp1661;
  assign tmp1661 = (tmp1658 & tmp1659) | (tmp1658 & tmp1660) | (tmp1659 & tmp1660);
  wire tmp1662;
  assign tmp1662 = 1'b1;
  wire tmp1663;
  assign tmp1663 = 1'b1;
  wire tmp1664;
  assign tmp1664 = 1'b1;
  wire tmp1665;
  assign tmp1665 = (tmp1662 & tmp1663) | (tmp1662 & tmp1664) | (tmp1663 & tmp1664);
  wire tmp1666;
  assign tmp1666 = 1'b0;
  wire tmp1667;
  assign tmp1667 = 1'b1;
  wire tmp1668;
  assign tmp1668 = 1'b0;
  wire tmp1669;
  assign tmp1669 = (tmp1666 & tmp1667) | (tmp1666 & tmp1668) | (tmp1667 & tmp1668);
  wire tmp1670;
  assign tmp1670 = (tmp1661 & tmp1665) | (tmp1661 & tmp1669) | (tmp1665 & tmp1669);
  wire tmp1671;
  assign tmp1671 = 1'b1;
  wire tmp1672;
  assign tmp1672 = 1'b1;
  wire tmp1673;
  assign tmp1673 = 1'b1;
  wire tmp1674;
  assign tmp1674 = (tmp1671 & tmp1672) | (tmp1671 & tmp1673) | (tmp1672 & tmp1673);
  wire tmp1675;
  assign tmp1675 = 1'b1;
  wire tmp1676;
  assign tmp1676 = ~pi5;
  wire tmp1677;
  assign tmp1677 = ~pi6;
  wire tmp1678;
  assign tmp1678 = (tmp1675 & tmp1676) | (tmp1675 & tmp1677) | (tmp1676 & tmp1677);
  wire tmp1679;
  assign tmp1679 = 1'b1;
  wire tmp1680;
  assign tmp1680 = ~pi6;
  wire tmp1681;
  assign tmp1681 = ~pi7;
  wire tmp1682;
  assign tmp1682 = (tmp1679 & tmp1680) | (tmp1679 & tmp1681) | (tmp1680 & tmp1681);
  wire tmp1683;
  assign tmp1683 = (tmp1674 & tmp1678) | (tmp1674 & tmp1682) | (tmp1678 & tmp1682);
  wire tmp1684;
  assign tmp1684 = 1'b0;
  wire tmp1685;
  assign tmp1685 = 1'b1;
  wire tmp1686;
  assign tmp1686 = 1'b0;
  wire tmp1687;
  assign tmp1687 = (tmp1684 & tmp1685) | (tmp1684 & tmp1686) | (tmp1685 & tmp1686);
  wire tmp1688;
  assign tmp1688 = 1'b1;
  wire tmp1689;
  assign tmp1689 = ~pi6;
  wire tmp1690;
  assign tmp1690 = ~pi7;
  wire tmp1691;
  assign tmp1691 = (tmp1688 & tmp1689) | (tmp1688 & tmp1690) | (tmp1689 & tmp1690);
  wire tmp1692;
  assign tmp1692 = 1'b0;
  wire tmp1693;
  assign tmp1693 = ~pi7;
  wire tmp1694;
  assign tmp1694 = 1'b0;
  wire tmp1695;
  assign tmp1695 = (tmp1692 & tmp1693) | (tmp1692 & tmp1694) | (tmp1693 & tmp1694);
  wire tmp1696;
  assign tmp1696 = (tmp1687 & tmp1691) | (tmp1687 & tmp1695) | (tmp1691 & tmp1695);
  wire tmp1697;
  assign tmp1697 = (tmp1670 & tmp1683) | (tmp1670 & tmp1696) | (tmp1683 & tmp1696);
  wire tmp1698;
  assign tmp1698 = (tmp1617 & tmp1657) | (tmp1617 & tmp1697) | (tmp1657 & tmp1697);
  wire tmp1699;
  assign tmp1699 = 1'b0;
  wire tmp1700;
  assign tmp1700 = 1'b0;
  wire tmp1701;
  assign tmp1701 = 1'b0;
  wire tmp1702;
  assign tmp1702 = (tmp1699 & tmp1700) | (tmp1699 & tmp1701) | (tmp1700 & tmp1701);
  wire tmp1703;
  assign tmp1703 = 1'b0;
  wire tmp1704;
  assign tmp1704 = 1'b1;
  wire tmp1705;
  assign tmp1705 = 1'b0;
  wire tmp1706;
  assign tmp1706 = (tmp1703 & tmp1704) | (tmp1703 & tmp1705) | (tmp1704 & tmp1705);
  wire tmp1707;
  assign tmp1707 = 1'b0;
  wire tmp1708;
  assign tmp1708 = 1'b0;
  wire tmp1709;
  assign tmp1709 = 1'b0;
  wire tmp1710;
  assign tmp1710 = (tmp1707 & tmp1708) | (tmp1707 & tmp1709) | (tmp1708 & tmp1709);
  wire tmp1711;
  assign tmp1711 = (tmp1702 & tmp1706) | (tmp1702 & tmp1710) | (tmp1706 & tmp1710);
  wire tmp1712;
  assign tmp1712 = 1'b0;
  wire tmp1713;
  assign tmp1713 = 1'b1;
  wire tmp1714;
  assign tmp1714 = 1'b0;
  wire tmp1715;
  assign tmp1715 = (tmp1712 & tmp1713) | (tmp1712 & tmp1714) | (tmp1713 & tmp1714);
  wire tmp1716;
  assign tmp1716 = 1'b1;
  wire tmp1717;
  assign tmp1717 = 1'b1;
  wire tmp1718;
  assign tmp1718 = 1'b1;
  wire tmp1719;
  assign tmp1719 = (tmp1716 & tmp1717) | (tmp1716 & tmp1718) | (tmp1717 & tmp1718);
  wire tmp1720;
  assign tmp1720 = 1'b0;
  wire tmp1721;
  assign tmp1721 = 1'b1;
  wire tmp1722;
  assign tmp1722 = 1'b0;
  wire tmp1723;
  assign tmp1723 = (tmp1720 & tmp1721) | (tmp1720 & tmp1722) | (tmp1721 & tmp1722);
  wire tmp1724;
  assign tmp1724 = (tmp1715 & tmp1719) | (tmp1715 & tmp1723) | (tmp1719 & tmp1723);
  wire tmp1725;
  assign tmp1725 = 1'b0;
  wire tmp1726;
  assign tmp1726 = 1'b0;
  wire tmp1727;
  assign tmp1727 = 1'b0;
  wire tmp1728;
  assign tmp1728 = (tmp1725 & tmp1726) | (tmp1725 & tmp1727) | (tmp1726 & tmp1727);
  wire tmp1729;
  assign tmp1729 = 1'b0;
  wire tmp1730;
  assign tmp1730 = 1'b1;
  wire tmp1731;
  assign tmp1731 = 1'b0;
  wire tmp1732;
  assign tmp1732 = (tmp1729 & tmp1730) | (tmp1729 & tmp1731) | (tmp1730 & tmp1731);
  wire tmp1733;
  assign tmp1733 = 1'b0;
  wire tmp1734;
  assign tmp1734 = 1'b0;
  wire tmp1735;
  assign tmp1735 = 1'b0;
  wire tmp1736;
  assign tmp1736 = (tmp1733 & tmp1734) | (tmp1733 & tmp1735) | (tmp1734 & tmp1735);
  wire tmp1737;
  assign tmp1737 = (tmp1728 & tmp1732) | (tmp1728 & tmp1736) | (tmp1732 & tmp1736);
  wire tmp1738;
  assign tmp1738 = (tmp1711 & tmp1724) | (tmp1711 & tmp1737) | (tmp1724 & tmp1737);
  wire tmp1739;
  assign tmp1739 = 1'b0;
  wire tmp1740;
  assign tmp1740 = 1'b1;
  wire tmp1741;
  assign tmp1741 = 1'b0;
  wire tmp1742;
  assign tmp1742 = (tmp1739 & tmp1740) | (tmp1739 & tmp1741) | (tmp1740 & tmp1741);
  wire tmp1743;
  assign tmp1743 = 1'b1;
  wire tmp1744;
  assign tmp1744 = 1'b1;
  wire tmp1745;
  assign tmp1745 = 1'b1;
  wire tmp1746;
  assign tmp1746 = (tmp1743 & tmp1744) | (tmp1743 & tmp1745) | (tmp1744 & tmp1745);
  wire tmp1747;
  assign tmp1747 = 1'b0;
  wire tmp1748;
  assign tmp1748 = 1'b1;
  wire tmp1749;
  assign tmp1749 = 1'b0;
  wire tmp1750;
  assign tmp1750 = (tmp1747 & tmp1748) | (tmp1747 & tmp1749) | (tmp1748 & tmp1749);
  wire tmp1751;
  assign tmp1751 = (tmp1742 & tmp1746) | (tmp1742 & tmp1750) | (tmp1746 & tmp1750);
  wire tmp1752;
  assign tmp1752 = 1'b1;
  wire tmp1753;
  assign tmp1753 = 1'b1;
  wire tmp1754;
  assign tmp1754 = 1'b1;
  wire tmp1755;
  assign tmp1755 = (tmp1752 & tmp1753) | (tmp1752 & tmp1754) | (tmp1753 & tmp1754);
  wire tmp1756;
  assign tmp1756 = 1'b1;
  wire tmp1757;
  assign tmp1757 = ~pi5;
  wire tmp1758;
  assign tmp1758 = ~pi6;
  wire tmp1759;
  assign tmp1759 = (tmp1756 & tmp1757) | (tmp1756 & tmp1758) | (tmp1757 & tmp1758);
  wire tmp1760;
  assign tmp1760 = 1'b1;
  wire tmp1761;
  assign tmp1761 = ~pi6;
  wire tmp1762;
  assign tmp1762 = ~pi7;
  wire tmp1763;
  assign tmp1763 = (tmp1760 & tmp1761) | (tmp1760 & tmp1762) | (tmp1761 & tmp1762);
  wire tmp1764;
  assign tmp1764 = (tmp1755 & tmp1759) | (tmp1755 & tmp1763) | (tmp1759 & tmp1763);
  wire tmp1765;
  assign tmp1765 = 1'b0;
  wire tmp1766;
  assign tmp1766 = 1'b1;
  wire tmp1767;
  assign tmp1767 = 1'b0;
  wire tmp1768;
  assign tmp1768 = (tmp1765 & tmp1766) | (tmp1765 & tmp1767) | (tmp1766 & tmp1767);
  wire tmp1769;
  assign tmp1769 = 1'b1;
  wire tmp1770;
  assign tmp1770 = ~pi6;
  wire tmp1771;
  assign tmp1771 = ~pi7;
  wire tmp1772;
  assign tmp1772 = (tmp1769 & tmp1770) | (tmp1769 & tmp1771) | (tmp1770 & tmp1771);
  wire tmp1773;
  assign tmp1773 = 1'b0;
  wire tmp1774;
  assign tmp1774 = ~pi7;
  wire tmp1775;
  assign tmp1775 = 1'b0;
  wire tmp1776;
  assign tmp1776 = (tmp1773 & tmp1774) | (tmp1773 & tmp1775) | (tmp1774 & tmp1775);
  wire tmp1777;
  assign tmp1777 = (tmp1768 & tmp1772) | (tmp1768 & tmp1776) | (tmp1772 & tmp1776);
  wire tmp1778;
  assign tmp1778 = (tmp1751 & tmp1764) | (tmp1751 & tmp1777) | (tmp1764 & tmp1777);
  wire tmp1779;
  assign tmp1779 = 1'b0;
  wire tmp1780;
  assign tmp1780 = 1'b0;
  wire tmp1781;
  assign tmp1781 = 1'b0;
  wire tmp1782;
  assign tmp1782 = (tmp1779 & tmp1780) | (tmp1779 & tmp1781) | (tmp1780 & tmp1781);
  wire tmp1783;
  assign tmp1783 = 1'b0;
  wire tmp1784;
  assign tmp1784 = 1'b1;
  wire tmp1785;
  assign tmp1785 = 1'b0;
  wire tmp1786;
  assign tmp1786 = (tmp1783 & tmp1784) | (tmp1783 & tmp1785) | (tmp1784 & tmp1785);
  wire tmp1787;
  assign tmp1787 = 1'b0;
  wire tmp1788;
  assign tmp1788 = 1'b0;
  wire tmp1789;
  assign tmp1789 = 1'b0;
  wire tmp1790;
  assign tmp1790 = (tmp1787 & tmp1788) | (tmp1787 & tmp1789) | (tmp1788 & tmp1789);
  wire tmp1791;
  assign tmp1791 = (tmp1782 & tmp1786) | (tmp1782 & tmp1790) | (tmp1786 & tmp1790);
  wire tmp1792;
  assign tmp1792 = 1'b0;
  wire tmp1793;
  assign tmp1793 = 1'b1;
  wire tmp1794;
  assign tmp1794 = 1'b0;
  wire tmp1795;
  assign tmp1795 = (tmp1792 & tmp1793) | (tmp1792 & tmp1794) | (tmp1793 & tmp1794);
  wire tmp1796;
  assign tmp1796 = 1'b1;
  wire tmp1797;
  assign tmp1797 = ~pi6;
  wire tmp1798;
  assign tmp1798 = ~pi7;
  wire tmp1799;
  assign tmp1799 = (tmp1796 & tmp1797) | (tmp1796 & tmp1798) | (tmp1797 & tmp1798);
  wire tmp1800;
  assign tmp1800 = 1'b0;
  wire tmp1801;
  assign tmp1801 = ~pi7;
  wire tmp1802;
  assign tmp1802 = 1'b0;
  wire tmp1803;
  assign tmp1803 = (tmp1800 & tmp1801) | (tmp1800 & tmp1802) | (tmp1801 & tmp1802);
  wire tmp1804;
  assign tmp1804 = (tmp1795 & tmp1799) | (tmp1795 & tmp1803) | (tmp1799 & tmp1803);
  wire tmp1805;
  assign tmp1805 = 1'b0;
  wire tmp1806;
  assign tmp1806 = 1'b0;
  wire tmp1807;
  assign tmp1807 = 1'b0;
  wire tmp1808;
  assign tmp1808 = (tmp1805 & tmp1806) | (tmp1805 & tmp1807) | (tmp1806 & tmp1807);
  wire tmp1809;
  assign tmp1809 = 1'b0;
  wire tmp1810;
  assign tmp1810 = ~pi7;
  wire tmp1811;
  assign tmp1811 = 1'b0;
  wire tmp1812;
  assign tmp1812 = (tmp1809 & tmp1810) | (tmp1809 & tmp1811) | (tmp1810 & tmp1811);
  wire tmp1813;
  assign tmp1813 = 1'b0;
  wire tmp1814;
  assign tmp1814 = 1'b0;
  wire tmp1815;
  assign tmp1815 = 1'b0;
  wire tmp1816;
  assign tmp1816 = (tmp1813 & tmp1814) | (tmp1813 & tmp1815) | (tmp1814 & tmp1815);
  wire tmp1817;
  assign tmp1817 = (tmp1808 & tmp1812) | (tmp1808 & tmp1816) | (tmp1812 & tmp1816);
  wire tmp1818;
  assign tmp1818 = (tmp1791 & tmp1804) | (tmp1791 & tmp1817) | (tmp1804 & tmp1817);
  wire tmp1819;
  assign tmp1819 = (tmp1738 & tmp1778) | (tmp1738 & tmp1818) | (tmp1778 & tmp1818);
  wire tmp1820;
  assign tmp1820 = (tmp1577 & tmp1698) | (tmp1577 & tmp1819) | (tmp1698 & tmp1819);
  wire tmp1821;
  assign tmp1821 = 1'b0;
  wire tmp1822;
  assign tmp1822 = 1'b0;
  wire tmp1823;
  assign tmp1823 = 1'b0;
  wire tmp1824;
  assign tmp1824 = (tmp1821 & tmp1822) | (tmp1821 & tmp1823) | (tmp1822 & tmp1823);
  wire tmp1825;
  assign tmp1825 = 1'b0;
  wire tmp1826;
  assign tmp1826 = 1'b0;
  wire tmp1827;
  assign tmp1827 = 1'b0;
  wire tmp1828;
  assign tmp1828 = (tmp1825 & tmp1826) | (tmp1825 & tmp1827) | (tmp1826 & tmp1827);
  wire tmp1829;
  assign tmp1829 = 1'b0;
  wire tmp1830;
  assign tmp1830 = 1'b0;
  wire tmp1831;
  assign tmp1831 = 1'b0;
  wire tmp1832;
  assign tmp1832 = (tmp1829 & tmp1830) | (tmp1829 & tmp1831) | (tmp1830 & tmp1831);
  wire tmp1833;
  assign tmp1833 = (tmp1824 & tmp1828) | (tmp1824 & tmp1832) | (tmp1828 & tmp1832);
  wire tmp1834;
  assign tmp1834 = 1'b0;
  wire tmp1835;
  assign tmp1835 = 1'b0;
  wire tmp1836;
  assign tmp1836 = 1'b0;
  wire tmp1837;
  assign tmp1837 = (tmp1834 & tmp1835) | (tmp1834 & tmp1836) | (tmp1835 & tmp1836);
  wire tmp1838;
  assign tmp1838 = 1'b0;
  wire tmp1839;
  assign tmp1839 = 1'b1;
  wire tmp1840;
  assign tmp1840 = 1'b0;
  wire tmp1841;
  assign tmp1841 = (tmp1838 & tmp1839) | (tmp1838 & tmp1840) | (tmp1839 & tmp1840);
  wire tmp1842;
  assign tmp1842 = 1'b0;
  wire tmp1843;
  assign tmp1843 = 1'b0;
  wire tmp1844;
  assign tmp1844 = 1'b0;
  wire tmp1845;
  assign tmp1845 = (tmp1842 & tmp1843) | (tmp1842 & tmp1844) | (tmp1843 & tmp1844);
  wire tmp1846;
  assign tmp1846 = (tmp1837 & tmp1841) | (tmp1837 & tmp1845) | (tmp1841 & tmp1845);
  wire tmp1847;
  assign tmp1847 = 1'b0;
  wire tmp1848;
  assign tmp1848 = 1'b0;
  wire tmp1849;
  assign tmp1849 = 1'b0;
  wire tmp1850;
  assign tmp1850 = (tmp1847 & tmp1848) | (tmp1847 & tmp1849) | (tmp1848 & tmp1849);
  wire tmp1851;
  assign tmp1851 = 1'b0;
  wire tmp1852;
  assign tmp1852 = 1'b0;
  wire tmp1853;
  assign tmp1853 = 1'b0;
  wire tmp1854;
  assign tmp1854 = (tmp1851 & tmp1852) | (tmp1851 & tmp1853) | (tmp1852 & tmp1853);
  wire tmp1855;
  assign tmp1855 = 1'b0;
  wire tmp1856;
  assign tmp1856 = 1'b0;
  wire tmp1857;
  assign tmp1857 = 1'b0;
  wire tmp1858;
  assign tmp1858 = (tmp1855 & tmp1856) | (tmp1855 & tmp1857) | (tmp1856 & tmp1857);
  wire tmp1859;
  assign tmp1859 = (tmp1850 & tmp1854) | (tmp1850 & tmp1858) | (tmp1854 & tmp1858);
  wire tmp1860;
  assign tmp1860 = (tmp1833 & tmp1846) | (tmp1833 & tmp1859) | (tmp1846 & tmp1859);
  wire tmp1861;
  assign tmp1861 = 1'b0;
  wire tmp1862;
  assign tmp1862 = 1'b0;
  wire tmp1863;
  assign tmp1863 = 1'b0;
  wire tmp1864;
  assign tmp1864 = (tmp1861 & tmp1862) | (tmp1861 & tmp1863) | (tmp1862 & tmp1863);
  wire tmp1865;
  assign tmp1865 = 1'b0;
  wire tmp1866;
  assign tmp1866 = 1'b1;
  wire tmp1867;
  assign tmp1867 = 1'b0;
  wire tmp1868;
  assign tmp1868 = (tmp1865 & tmp1866) | (tmp1865 & tmp1867) | (tmp1866 & tmp1867);
  wire tmp1869;
  assign tmp1869 = 1'b0;
  wire tmp1870;
  assign tmp1870 = 1'b0;
  wire tmp1871;
  assign tmp1871 = 1'b0;
  wire tmp1872;
  assign tmp1872 = (tmp1869 & tmp1870) | (tmp1869 & tmp1871) | (tmp1870 & tmp1871);
  wire tmp1873;
  assign tmp1873 = (tmp1864 & tmp1868) | (tmp1864 & tmp1872) | (tmp1868 & tmp1872);
  wire tmp1874;
  assign tmp1874 = 1'b0;
  wire tmp1875;
  assign tmp1875 = 1'b1;
  wire tmp1876;
  assign tmp1876 = 1'b0;
  wire tmp1877;
  assign tmp1877 = (tmp1874 & tmp1875) | (tmp1874 & tmp1876) | (tmp1875 & tmp1876);
  wire tmp1878;
  assign tmp1878 = 1'b1;
  wire tmp1879;
  assign tmp1879 = 1'b1;
  wire tmp1880;
  assign tmp1880 = 1'b1;
  wire tmp1881;
  assign tmp1881 = (tmp1878 & tmp1879) | (tmp1878 & tmp1880) | (tmp1879 & tmp1880);
  wire tmp1882;
  assign tmp1882 = 1'b0;
  wire tmp1883;
  assign tmp1883 = 1'b1;
  wire tmp1884;
  assign tmp1884 = 1'b0;
  wire tmp1885;
  assign tmp1885 = (tmp1882 & tmp1883) | (tmp1882 & tmp1884) | (tmp1883 & tmp1884);
  wire tmp1886;
  assign tmp1886 = (tmp1877 & tmp1881) | (tmp1877 & tmp1885) | (tmp1881 & tmp1885);
  wire tmp1887;
  assign tmp1887 = 1'b0;
  wire tmp1888;
  assign tmp1888 = 1'b0;
  wire tmp1889;
  assign tmp1889 = 1'b0;
  wire tmp1890;
  assign tmp1890 = (tmp1887 & tmp1888) | (tmp1887 & tmp1889) | (tmp1888 & tmp1889);
  wire tmp1891;
  assign tmp1891 = 1'b0;
  wire tmp1892;
  assign tmp1892 = 1'b1;
  wire tmp1893;
  assign tmp1893 = 1'b0;
  wire tmp1894;
  assign tmp1894 = (tmp1891 & tmp1892) | (tmp1891 & tmp1893) | (tmp1892 & tmp1893);
  wire tmp1895;
  assign tmp1895 = 1'b0;
  wire tmp1896;
  assign tmp1896 = 1'b0;
  wire tmp1897;
  assign tmp1897 = 1'b0;
  wire tmp1898;
  assign tmp1898 = (tmp1895 & tmp1896) | (tmp1895 & tmp1897) | (tmp1896 & tmp1897);
  wire tmp1899;
  assign tmp1899 = (tmp1890 & tmp1894) | (tmp1890 & tmp1898) | (tmp1894 & tmp1898);
  wire tmp1900;
  assign tmp1900 = (tmp1873 & tmp1886) | (tmp1873 & tmp1899) | (tmp1886 & tmp1899);
  wire tmp1901;
  assign tmp1901 = 1'b0;
  wire tmp1902;
  assign tmp1902 = 1'b0;
  wire tmp1903;
  assign tmp1903 = 1'b0;
  wire tmp1904;
  assign tmp1904 = (tmp1901 & tmp1902) | (tmp1901 & tmp1903) | (tmp1902 & tmp1903);
  wire tmp1905;
  assign tmp1905 = 1'b0;
  wire tmp1906;
  assign tmp1906 = 1'b0;
  wire tmp1907;
  assign tmp1907 = 1'b0;
  wire tmp1908;
  assign tmp1908 = (tmp1905 & tmp1906) | (tmp1905 & tmp1907) | (tmp1906 & tmp1907);
  wire tmp1909;
  assign tmp1909 = 1'b0;
  wire tmp1910;
  assign tmp1910 = 1'b0;
  wire tmp1911;
  assign tmp1911 = 1'b0;
  wire tmp1912;
  assign tmp1912 = (tmp1909 & tmp1910) | (tmp1909 & tmp1911) | (tmp1910 & tmp1911);
  wire tmp1913;
  assign tmp1913 = (tmp1904 & tmp1908) | (tmp1904 & tmp1912) | (tmp1908 & tmp1912);
  wire tmp1914;
  assign tmp1914 = 1'b0;
  wire tmp1915;
  assign tmp1915 = 1'b0;
  wire tmp1916;
  assign tmp1916 = 1'b0;
  wire tmp1917;
  assign tmp1917 = (tmp1914 & tmp1915) | (tmp1914 & tmp1916) | (tmp1915 & tmp1916);
  wire tmp1918;
  assign tmp1918 = 1'b0;
  wire tmp1919;
  assign tmp1919 = 1'b1;
  wire tmp1920;
  assign tmp1920 = 1'b0;
  wire tmp1921;
  assign tmp1921 = (tmp1918 & tmp1919) | (tmp1918 & tmp1920) | (tmp1919 & tmp1920);
  wire tmp1922;
  assign tmp1922 = 1'b0;
  wire tmp1923;
  assign tmp1923 = 1'b0;
  wire tmp1924;
  assign tmp1924 = 1'b0;
  wire tmp1925;
  assign tmp1925 = (tmp1922 & tmp1923) | (tmp1922 & tmp1924) | (tmp1923 & tmp1924);
  wire tmp1926;
  assign tmp1926 = (tmp1917 & tmp1921) | (tmp1917 & tmp1925) | (tmp1921 & tmp1925);
  wire tmp1927;
  assign tmp1927 = 1'b0;
  wire tmp1928;
  assign tmp1928 = 1'b0;
  wire tmp1929;
  assign tmp1929 = 1'b0;
  wire tmp1930;
  assign tmp1930 = (tmp1927 & tmp1928) | (tmp1927 & tmp1929) | (tmp1928 & tmp1929);
  wire tmp1931;
  assign tmp1931 = 1'b0;
  wire tmp1932;
  assign tmp1932 = 1'b0;
  wire tmp1933;
  assign tmp1933 = 1'b0;
  wire tmp1934;
  assign tmp1934 = (tmp1931 & tmp1932) | (tmp1931 & tmp1933) | (tmp1932 & tmp1933);
  wire tmp1935;
  assign tmp1935 = 1'b0;
  wire tmp1936;
  assign tmp1936 = 1'b0;
  wire tmp1937;
  assign tmp1937 = 1'b0;
  wire tmp1938;
  assign tmp1938 = (tmp1935 & tmp1936) | (tmp1935 & tmp1937) | (tmp1936 & tmp1937);
  wire tmp1939;
  assign tmp1939 = (tmp1930 & tmp1934) | (tmp1930 & tmp1938) | (tmp1934 & tmp1938);
  wire tmp1940;
  assign tmp1940 = (tmp1913 & tmp1926) | (tmp1913 & tmp1939) | (tmp1926 & tmp1939);
  wire tmp1941;
  assign tmp1941 = (tmp1860 & tmp1900) | (tmp1860 & tmp1940) | (tmp1900 & tmp1940);
  wire tmp1942;
  assign tmp1942 = 1'b0;
  wire tmp1943;
  assign tmp1943 = 1'b0;
  wire tmp1944;
  assign tmp1944 = 1'b0;
  wire tmp1945;
  assign tmp1945 = (tmp1942 & tmp1943) | (tmp1942 & tmp1944) | (tmp1943 & tmp1944);
  wire tmp1946;
  assign tmp1946 = 1'b0;
  wire tmp1947;
  assign tmp1947 = 1'b1;
  wire tmp1948;
  assign tmp1948 = 1'b0;
  wire tmp1949;
  assign tmp1949 = (tmp1946 & tmp1947) | (tmp1946 & tmp1948) | (tmp1947 & tmp1948);
  wire tmp1950;
  assign tmp1950 = 1'b0;
  wire tmp1951;
  assign tmp1951 = 1'b0;
  wire tmp1952;
  assign tmp1952 = 1'b0;
  wire tmp1953;
  assign tmp1953 = (tmp1950 & tmp1951) | (tmp1950 & tmp1952) | (tmp1951 & tmp1952);
  wire tmp1954;
  assign tmp1954 = (tmp1945 & tmp1949) | (tmp1945 & tmp1953) | (tmp1949 & tmp1953);
  wire tmp1955;
  assign tmp1955 = 1'b0;
  wire tmp1956;
  assign tmp1956 = 1'b1;
  wire tmp1957;
  assign tmp1957 = 1'b0;
  wire tmp1958;
  assign tmp1958 = (tmp1955 & tmp1956) | (tmp1955 & tmp1957) | (tmp1956 & tmp1957);
  wire tmp1959;
  assign tmp1959 = 1'b1;
  wire tmp1960;
  assign tmp1960 = 1'b1;
  wire tmp1961;
  assign tmp1961 = 1'b1;
  wire tmp1962;
  assign tmp1962 = (tmp1959 & tmp1960) | (tmp1959 & tmp1961) | (tmp1960 & tmp1961);
  wire tmp1963;
  assign tmp1963 = 1'b0;
  wire tmp1964;
  assign tmp1964 = 1'b1;
  wire tmp1965;
  assign tmp1965 = 1'b0;
  wire tmp1966;
  assign tmp1966 = (tmp1963 & tmp1964) | (tmp1963 & tmp1965) | (tmp1964 & tmp1965);
  wire tmp1967;
  assign tmp1967 = (tmp1958 & tmp1962) | (tmp1958 & tmp1966) | (tmp1962 & tmp1966);
  wire tmp1968;
  assign tmp1968 = 1'b0;
  wire tmp1969;
  assign tmp1969 = 1'b0;
  wire tmp1970;
  assign tmp1970 = 1'b0;
  wire tmp1971;
  assign tmp1971 = (tmp1968 & tmp1969) | (tmp1968 & tmp1970) | (tmp1969 & tmp1970);
  wire tmp1972;
  assign tmp1972 = 1'b0;
  wire tmp1973;
  assign tmp1973 = 1'b1;
  wire tmp1974;
  assign tmp1974 = 1'b0;
  wire tmp1975;
  assign tmp1975 = (tmp1972 & tmp1973) | (tmp1972 & tmp1974) | (tmp1973 & tmp1974);
  wire tmp1976;
  assign tmp1976 = 1'b0;
  wire tmp1977;
  assign tmp1977 = 1'b0;
  wire tmp1978;
  assign tmp1978 = 1'b0;
  wire tmp1979;
  assign tmp1979 = (tmp1976 & tmp1977) | (tmp1976 & tmp1978) | (tmp1977 & tmp1978);
  wire tmp1980;
  assign tmp1980 = (tmp1971 & tmp1975) | (tmp1971 & tmp1979) | (tmp1975 & tmp1979);
  wire tmp1981;
  assign tmp1981 = (tmp1954 & tmp1967) | (tmp1954 & tmp1980) | (tmp1967 & tmp1980);
  wire tmp1982;
  assign tmp1982 = 1'b0;
  wire tmp1983;
  assign tmp1983 = 1'b1;
  wire tmp1984;
  assign tmp1984 = 1'b0;
  wire tmp1985;
  assign tmp1985 = (tmp1982 & tmp1983) | (tmp1982 & tmp1984) | (tmp1983 & tmp1984);
  wire tmp1986;
  assign tmp1986 = 1'b1;
  wire tmp1987;
  assign tmp1987 = 1'b1;
  wire tmp1988;
  assign tmp1988 = 1'b1;
  wire tmp1989;
  assign tmp1989 = (tmp1986 & tmp1987) | (tmp1986 & tmp1988) | (tmp1987 & tmp1988);
  wire tmp1990;
  assign tmp1990 = 1'b0;
  wire tmp1991;
  assign tmp1991 = 1'b1;
  wire tmp1992;
  assign tmp1992 = 1'b0;
  wire tmp1993;
  assign tmp1993 = (tmp1990 & tmp1991) | (tmp1990 & tmp1992) | (tmp1991 & tmp1992);
  wire tmp1994;
  assign tmp1994 = (tmp1985 & tmp1989) | (tmp1985 & tmp1993) | (tmp1989 & tmp1993);
  wire tmp1995;
  assign tmp1995 = 1'b1;
  wire tmp1996;
  assign tmp1996 = 1'b1;
  wire tmp1997;
  assign tmp1997 = 1'b1;
  wire tmp1998;
  assign tmp1998 = (tmp1995 & tmp1996) | (tmp1995 & tmp1997) | (tmp1996 & tmp1997);
  wire tmp1999;
  assign tmp1999 = 1'b1;
  wire tmp2000;
  assign tmp2000 = ~pi5;
  wire tmp2001;
  assign tmp2001 = ~pi6;
  wire tmp2002;
  assign tmp2002 = (tmp1999 & tmp2000) | (tmp1999 & tmp2001) | (tmp2000 & tmp2001);
  wire tmp2003;
  assign tmp2003 = 1'b1;
  wire tmp2004;
  assign tmp2004 = ~pi6;
  wire tmp2005;
  assign tmp2005 = ~pi7;
  wire tmp2006;
  assign tmp2006 = (tmp2003 & tmp2004) | (tmp2003 & tmp2005) | (tmp2004 & tmp2005);
  wire tmp2007;
  assign tmp2007 = (tmp1998 & tmp2002) | (tmp1998 & tmp2006) | (tmp2002 & tmp2006);
  wire tmp2008;
  assign tmp2008 = 1'b0;
  wire tmp2009;
  assign tmp2009 = 1'b1;
  wire tmp2010;
  assign tmp2010 = 1'b0;
  wire tmp2011;
  assign tmp2011 = (tmp2008 & tmp2009) | (tmp2008 & tmp2010) | (tmp2009 & tmp2010);
  wire tmp2012;
  assign tmp2012 = 1'b1;
  wire tmp2013;
  assign tmp2013 = ~pi6;
  wire tmp2014;
  assign tmp2014 = ~pi7;
  wire tmp2015;
  assign tmp2015 = (tmp2012 & tmp2013) | (tmp2012 & tmp2014) | (tmp2013 & tmp2014);
  wire tmp2016;
  assign tmp2016 = 1'b0;
  wire tmp2017;
  assign tmp2017 = ~pi7;
  wire tmp2018;
  assign tmp2018 = 1'b0;
  wire tmp2019;
  assign tmp2019 = (tmp2016 & tmp2017) | (tmp2016 & tmp2018) | (tmp2017 & tmp2018);
  wire tmp2020;
  assign tmp2020 = (tmp2011 & tmp2015) | (tmp2011 & tmp2019) | (tmp2015 & tmp2019);
  wire tmp2021;
  assign tmp2021 = (tmp1994 & tmp2007) | (tmp1994 & tmp2020) | (tmp2007 & tmp2020);
  wire tmp2022;
  assign tmp2022 = 1'b0;
  wire tmp2023;
  assign tmp2023 = 1'b0;
  wire tmp2024;
  assign tmp2024 = 1'b0;
  wire tmp2025;
  assign tmp2025 = (tmp2022 & tmp2023) | (tmp2022 & tmp2024) | (tmp2023 & tmp2024);
  wire tmp2026;
  assign tmp2026 = 1'b0;
  wire tmp2027;
  assign tmp2027 = 1'b1;
  wire tmp2028;
  assign tmp2028 = 1'b0;
  wire tmp2029;
  assign tmp2029 = (tmp2026 & tmp2027) | (tmp2026 & tmp2028) | (tmp2027 & tmp2028);
  wire tmp2030;
  assign tmp2030 = 1'b0;
  wire tmp2031;
  assign tmp2031 = 1'b0;
  wire tmp2032;
  assign tmp2032 = 1'b0;
  wire tmp2033;
  assign tmp2033 = (tmp2030 & tmp2031) | (tmp2030 & tmp2032) | (tmp2031 & tmp2032);
  wire tmp2034;
  assign tmp2034 = (tmp2025 & tmp2029) | (tmp2025 & tmp2033) | (tmp2029 & tmp2033);
  wire tmp2035;
  assign tmp2035 = 1'b0;
  wire tmp2036;
  assign tmp2036 = 1'b1;
  wire tmp2037;
  assign tmp2037 = 1'b0;
  wire tmp2038;
  assign tmp2038 = (tmp2035 & tmp2036) | (tmp2035 & tmp2037) | (tmp2036 & tmp2037);
  wire tmp2039;
  assign tmp2039 = 1'b1;
  wire tmp2040;
  assign tmp2040 = ~pi6;
  wire tmp2041;
  assign tmp2041 = ~pi7;
  wire tmp2042;
  assign tmp2042 = (tmp2039 & tmp2040) | (tmp2039 & tmp2041) | (tmp2040 & tmp2041);
  wire tmp2043;
  assign tmp2043 = 1'b0;
  wire tmp2044;
  assign tmp2044 = ~pi7;
  wire tmp2045;
  assign tmp2045 = 1'b0;
  wire tmp2046;
  assign tmp2046 = (tmp2043 & tmp2044) | (tmp2043 & tmp2045) | (tmp2044 & tmp2045);
  wire tmp2047;
  assign tmp2047 = (tmp2038 & tmp2042) | (tmp2038 & tmp2046) | (tmp2042 & tmp2046);
  wire tmp2048;
  assign tmp2048 = 1'b0;
  wire tmp2049;
  assign tmp2049 = 1'b0;
  wire tmp2050;
  assign tmp2050 = 1'b0;
  wire tmp2051;
  assign tmp2051 = (tmp2048 & tmp2049) | (tmp2048 & tmp2050) | (tmp2049 & tmp2050);
  wire tmp2052;
  assign tmp2052 = 1'b0;
  wire tmp2053;
  assign tmp2053 = ~pi7;
  wire tmp2054;
  assign tmp2054 = 1'b0;
  wire tmp2055;
  assign tmp2055 = (tmp2052 & tmp2053) | (tmp2052 & tmp2054) | (tmp2053 & tmp2054);
  wire tmp2056;
  assign tmp2056 = 1'b0;
  wire tmp2057;
  assign tmp2057 = 1'b0;
  wire tmp2058;
  assign tmp2058 = 1'b0;
  wire tmp2059;
  assign tmp2059 = (tmp2056 & tmp2057) | (tmp2056 & tmp2058) | (tmp2057 & tmp2058);
  wire tmp2060;
  assign tmp2060 = (tmp2051 & tmp2055) | (tmp2051 & tmp2059) | (tmp2055 & tmp2059);
  wire tmp2061;
  assign tmp2061 = (tmp2034 & tmp2047) | (tmp2034 & tmp2060) | (tmp2047 & tmp2060);
  wire tmp2062;
  assign tmp2062 = (tmp1981 & tmp2021) | (tmp1981 & tmp2061) | (tmp2021 & tmp2061);
  wire tmp2063;
  assign tmp2063 = 1'b0;
  wire tmp2064;
  assign tmp2064 = 1'b0;
  wire tmp2065;
  assign tmp2065 = 1'b0;
  wire tmp2066;
  assign tmp2066 = (tmp2063 & tmp2064) | (tmp2063 & tmp2065) | (tmp2064 & tmp2065);
  wire tmp2067;
  assign tmp2067 = 1'b0;
  wire tmp2068;
  assign tmp2068 = 1'b0;
  wire tmp2069;
  assign tmp2069 = 1'b0;
  wire tmp2070;
  assign tmp2070 = (tmp2067 & tmp2068) | (tmp2067 & tmp2069) | (tmp2068 & tmp2069);
  wire tmp2071;
  assign tmp2071 = 1'b0;
  wire tmp2072;
  assign tmp2072 = 1'b0;
  wire tmp2073;
  assign tmp2073 = 1'b0;
  wire tmp2074;
  assign tmp2074 = (tmp2071 & tmp2072) | (tmp2071 & tmp2073) | (tmp2072 & tmp2073);
  wire tmp2075;
  assign tmp2075 = (tmp2066 & tmp2070) | (tmp2066 & tmp2074) | (tmp2070 & tmp2074);
  wire tmp2076;
  assign tmp2076 = 1'b0;
  wire tmp2077;
  assign tmp2077 = 1'b0;
  wire tmp2078;
  assign tmp2078 = 1'b0;
  wire tmp2079;
  assign tmp2079 = (tmp2076 & tmp2077) | (tmp2076 & tmp2078) | (tmp2077 & tmp2078);
  wire tmp2080;
  assign tmp2080 = 1'b0;
  wire tmp2081;
  assign tmp2081 = 1'b1;
  wire tmp2082;
  assign tmp2082 = 1'b0;
  wire tmp2083;
  assign tmp2083 = (tmp2080 & tmp2081) | (tmp2080 & tmp2082) | (tmp2081 & tmp2082);
  wire tmp2084;
  assign tmp2084 = 1'b0;
  wire tmp2085;
  assign tmp2085 = 1'b0;
  wire tmp2086;
  assign tmp2086 = 1'b0;
  wire tmp2087;
  assign tmp2087 = (tmp2084 & tmp2085) | (tmp2084 & tmp2086) | (tmp2085 & tmp2086);
  wire tmp2088;
  assign tmp2088 = (tmp2079 & tmp2083) | (tmp2079 & tmp2087) | (tmp2083 & tmp2087);
  wire tmp2089;
  assign tmp2089 = 1'b0;
  wire tmp2090;
  assign tmp2090 = 1'b0;
  wire tmp2091;
  assign tmp2091 = 1'b0;
  wire tmp2092;
  assign tmp2092 = (tmp2089 & tmp2090) | (tmp2089 & tmp2091) | (tmp2090 & tmp2091);
  wire tmp2093;
  assign tmp2093 = 1'b0;
  wire tmp2094;
  assign tmp2094 = 1'b0;
  wire tmp2095;
  assign tmp2095 = 1'b0;
  wire tmp2096;
  assign tmp2096 = (tmp2093 & tmp2094) | (tmp2093 & tmp2095) | (tmp2094 & tmp2095);
  wire tmp2097;
  assign tmp2097 = 1'b0;
  wire tmp2098;
  assign tmp2098 = 1'b0;
  wire tmp2099;
  assign tmp2099 = 1'b0;
  wire tmp2100;
  assign tmp2100 = (tmp2097 & tmp2098) | (tmp2097 & tmp2099) | (tmp2098 & tmp2099);
  wire tmp2101;
  assign tmp2101 = (tmp2092 & tmp2096) | (tmp2092 & tmp2100) | (tmp2096 & tmp2100);
  wire tmp2102;
  assign tmp2102 = (tmp2075 & tmp2088) | (tmp2075 & tmp2101) | (tmp2088 & tmp2101);
  wire tmp2103;
  assign tmp2103 = 1'b0;
  wire tmp2104;
  assign tmp2104 = 1'b0;
  wire tmp2105;
  assign tmp2105 = 1'b0;
  wire tmp2106;
  assign tmp2106 = (tmp2103 & tmp2104) | (tmp2103 & tmp2105) | (tmp2104 & tmp2105);
  wire tmp2107;
  assign tmp2107 = 1'b0;
  wire tmp2108;
  assign tmp2108 = 1'b1;
  wire tmp2109;
  assign tmp2109 = 1'b0;
  wire tmp2110;
  assign tmp2110 = (tmp2107 & tmp2108) | (tmp2107 & tmp2109) | (tmp2108 & tmp2109);
  wire tmp2111;
  assign tmp2111 = 1'b0;
  wire tmp2112;
  assign tmp2112 = 1'b0;
  wire tmp2113;
  assign tmp2113 = 1'b0;
  wire tmp2114;
  assign tmp2114 = (tmp2111 & tmp2112) | (tmp2111 & tmp2113) | (tmp2112 & tmp2113);
  wire tmp2115;
  assign tmp2115 = (tmp2106 & tmp2110) | (tmp2106 & tmp2114) | (tmp2110 & tmp2114);
  wire tmp2116;
  assign tmp2116 = 1'b0;
  wire tmp2117;
  assign tmp2117 = 1'b1;
  wire tmp2118;
  assign tmp2118 = 1'b0;
  wire tmp2119;
  assign tmp2119 = (tmp2116 & tmp2117) | (tmp2116 & tmp2118) | (tmp2117 & tmp2118);
  wire tmp2120;
  assign tmp2120 = 1'b1;
  wire tmp2121;
  assign tmp2121 = ~pi6;
  wire tmp2122;
  assign tmp2122 = ~pi7;
  wire tmp2123;
  assign tmp2123 = (tmp2120 & tmp2121) | (tmp2120 & tmp2122) | (tmp2121 & tmp2122);
  wire tmp2124;
  assign tmp2124 = 1'b0;
  wire tmp2125;
  assign tmp2125 = ~pi7;
  wire tmp2126;
  assign tmp2126 = 1'b0;
  wire tmp2127;
  assign tmp2127 = (tmp2124 & tmp2125) | (tmp2124 & tmp2126) | (tmp2125 & tmp2126);
  wire tmp2128;
  assign tmp2128 = (tmp2119 & tmp2123) | (tmp2119 & tmp2127) | (tmp2123 & tmp2127);
  wire tmp2129;
  assign tmp2129 = 1'b0;
  wire tmp2130;
  assign tmp2130 = 1'b0;
  wire tmp2131;
  assign tmp2131 = 1'b0;
  wire tmp2132;
  assign tmp2132 = (tmp2129 & tmp2130) | (tmp2129 & tmp2131) | (tmp2130 & tmp2131);
  wire tmp2133;
  assign tmp2133 = 1'b0;
  wire tmp2134;
  assign tmp2134 = ~pi7;
  wire tmp2135;
  assign tmp2135 = 1'b0;
  wire tmp2136;
  assign tmp2136 = (tmp2133 & tmp2134) | (tmp2133 & tmp2135) | (tmp2134 & tmp2135);
  wire tmp2137;
  assign tmp2137 = 1'b0;
  wire tmp2138;
  assign tmp2138 = 1'b0;
  wire tmp2139;
  assign tmp2139 = 1'b0;
  wire tmp2140;
  assign tmp2140 = (tmp2137 & tmp2138) | (tmp2137 & tmp2139) | (tmp2138 & tmp2139);
  wire tmp2141;
  assign tmp2141 = (tmp2132 & tmp2136) | (tmp2132 & tmp2140) | (tmp2136 & tmp2140);
  wire tmp2142;
  assign tmp2142 = (tmp2115 & tmp2128) | (tmp2115 & tmp2141) | (tmp2128 & tmp2141);
  wire tmp2143;
  assign tmp2143 = 1'b0;
  wire tmp2144;
  assign tmp2144 = 1'b0;
  wire tmp2145;
  assign tmp2145 = 1'b0;
  wire tmp2146;
  assign tmp2146 = (tmp2143 & tmp2144) | (tmp2143 & tmp2145) | (tmp2144 & tmp2145);
  wire tmp2147;
  assign tmp2147 = 1'b0;
  wire tmp2148;
  assign tmp2148 = 1'b0;
  wire tmp2149;
  assign tmp2149 = 1'b0;
  wire tmp2150;
  assign tmp2150 = (tmp2147 & tmp2148) | (tmp2147 & tmp2149) | (tmp2148 & tmp2149);
  wire tmp2151;
  assign tmp2151 = 1'b0;
  wire tmp2152;
  assign tmp2152 = 1'b0;
  wire tmp2153;
  assign tmp2153 = 1'b0;
  wire tmp2154;
  assign tmp2154 = (tmp2151 & tmp2152) | (tmp2151 & tmp2153) | (tmp2152 & tmp2153);
  wire tmp2155;
  assign tmp2155 = (tmp2146 & tmp2150) | (tmp2146 & tmp2154) | (tmp2150 & tmp2154);
  wire tmp2156;
  assign tmp2156 = 1'b0;
  wire tmp2157;
  assign tmp2157 = 1'b0;
  wire tmp2158;
  assign tmp2158 = 1'b0;
  wire tmp2159;
  assign tmp2159 = (tmp2156 & tmp2157) | (tmp2156 & tmp2158) | (tmp2157 & tmp2158);
  wire tmp2160;
  assign tmp2160 = 1'b0;
  wire tmp2161;
  assign tmp2161 = ~pi7;
  wire tmp2162;
  assign tmp2162 = 1'b0;
  wire tmp2163;
  assign tmp2163 = (tmp2160 & tmp2161) | (tmp2160 & tmp2162) | (tmp2161 & tmp2162);
  wire tmp2164;
  assign tmp2164 = 1'b0;
  wire tmp2165;
  assign tmp2165 = 1'b0;
  wire tmp2166;
  assign tmp2166 = 1'b0;
  wire tmp2167;
  assign tmp2167 = (tmp2164 & tmp2165) | (tmp2164 & tmp2166) | (tmp2165 & tmp2166);
  wire tmp2168;
  assign tmp2168 = (tmp2159 & tmp2163) | (tmp2159 & tmp2167) | (tmp2163 & tmp2167);
  wire tmp2169;
  assign tmp2169 = 1'b0;
  wire tmp2170;
  assign tmp2170 = 1'b0;
  wire tmp2171;
  assign tmp2171 = 1'b0;
  wire tmp2172;
  assign tmp2172 = (tmp2169 & tmp2170) | (tmp2169 & tmp2171) | (tmp2170 & tmp2171);
  wire tmp2173;
  assign tmp2173 = 1'b0;
  wire tmp2174;
  assign tmp2174 = 1'b0;
  wire tmp2175;
  assign tmp2175 = 1'b0;
  wire tmp2176;
  assign tmp2176 = (tmp2173 & tmp2174) | (tmp2173 & tmp2175) | (tmp2174 & tmp2175);
  wire tmp2177;
  assign tmp2177 = 1'b0;
  wire tmp2178;
  assign tmp2178 = 1'b0;
  wire tmp2179;
  assign tmp2179 = 1'b0;
  wire tmp2180;
  assign tmp2180 = (tmp2177 & tmp2178) | (tmp2177 & tmp2179) | (tmp2178 & tmp2179);
  wire tmp2181;
  assign tmp2181 = (tmp2172 & tmp2176) | (tmp2172 & tmp2180) | (tmp2176 & tmp2180);
  wire tmp2182;
  assign tmp2182 = (tmp2155 & tmp2168) | (tmp2155 & tmp2181) | (tmp2168 & tmp2181);
  wire tmp2183;
  assign tmp2183 = (tmp2102 & tmp2142) | (tmp2102 & tmp2182) | (tmp2142 & tmp2182);
  wire tmp2184;
  assign tmp2184 = (tmp1941 & tmp2062) | (tmp1941 & tmp2183) | (tmp2062 & tmp2183);
  wire tmp2185;
  assign tmp2185 = (tmp1456 & tmp1820) | (tmp1456 & tmp2184) | (tmp1820 & tmp2184);
  wire tmp2186;
  assign tmp2186 = 1'b0;
  wire tmp2187;
  assign tmp2187 = 1'b0;
  wire tmp2188;
  assign tmp2188 = 1'b0;
  wire tmp2189;
  assign tmp2189 = (tmp2186 & tmp2187) | (tmp2186 & tmp2188) | (tmp2187 & tmp2188);
  wire tmp2190;
  assign tmp2190 = 1'b0;
  wire tmp2191;
  assign tmp2191 = 1'b0;
  wire tmp2192;
  assign tmp2192 = 1'b0;
  wire tmp2193;
  assign tmp2193 = (tmp2190 & tmp2191) | (tmp2190 & tmp2192) | (tmp2191 & tmp2192);
  wire tmp2194;
  assign tmp2194 = 1'b0;
  wire tmp2195;
  assign tmp2195 = 1'b0;
  wire tmp2196;
  assign tmp2196 = 1'b0;
  wire tmp2197;
  assign tmp2197 = (tmp2194 & tmp2195) | (tmp2194 & tmp2196) | (tmp2195 & tmp2196);
  wire tmp2198;
  assign tmp2198 = (tmp2189 & tmp2193) | (tmp2189 & tmp2197) | (tmp2193 & tmp2197);
  wire tmp2199;
  assign tmp2199 = 1'b0;
  wire tmp2200;
  assign tmp2200 = 1'b0;
  wire tmp2201;
  assign tmp2201 = 1'b0;
  wire tmp2202;
  assign tmp2202 = (tmp2199 & tmp2200) | (tmp2199 & tmp2201) | (tmp2200 & tmp2201);
  wire tmp2203;
  assign tmp2203 = 1'b0;
  wire tmp2204;
  assign tmp2204 = 1'b0;
  wire tmp2205;
  assign tmp2205 = 1'b0;
  wire tmp2206;
  assign tmp2206 = (tmp2203 & tmp2204) | (tmp2203 & tmp2205) | (tmp2204 & tmp2205);
  wire tmp2207;
  assign tmp2207 = 1'b0;
  wire tmp2208;
  assign tmp2208 = 1'b0;
  wire tmp2209;
  assign tmp2209 = 1'b0;
  wire tmp2210;
  assign tmp2210 = (tmp2207 & tmp2208) | (tmp2207 & tmp2209) | (tmp2208 & tmp2209);
  wire tmp2211;
  assign tmp2211 = (tmp2202 & tmp2206) | (tmp2202 & tmp2210) | (tmp2206 & tmp2210);
  wire tmp2212;
  assign tmp2212 = 1'b0;
  wire tmp2213;
  assign tmp2213 = 1'b0;
  wire tmp2214;
  assign tmp2214 = 1'b0;
  wire tmp2215;
  assign tmp2215 = (tmp2212 & tmp2213) | (tmp2212 & tmp2214) | (tmp2213 & tmp2214);
  wire tmp2216;
  assign tmp2216 = 1'b0;
  wire tmp2217;
  assign tmp2217 = 1'b0;
  wire tmp2218;
  assign tmp2218 = 1'b0;
  wire tmp2219;
  assign tmp2219 = (tmp2216 & tmp2217) | (tmp2216 & tmp2218) | (tmp2217 & tmp2218);
  wire tmp2220;
  assign tmp2220 = 1'b0;
  wire tmp2221;
  assign tmp2221 = 1'b0;
  wire tmp2222;
  assign tmp2222 = 1'b0;
  wire tmp2223;
  assign tmp2223 = (tmp2220 & tmp2221) | (tmp2220 & tmp2222) | (tmp2221 & tmp2222);
  wire tmp2224;
  assign tmp2224 = (tmp2215 & tmp2219) | (tmp2215 & tmp2223) | (tmp2219 & tmp2223);
  wire tmp2225;
  assign tmp2225 = (tmp2198 & tmp2211) | (tmp2198 & tmp2224) | (tmp2211 & tmp2224);
  wire tmp2226;
  assign tmp2226 = 1'b0;
  wire tmp2227;
  assign tmp2227 = 1'b0;
  wire tmp2228;
  assign tmp2228 = 1'b0;
  wire tmp2229;
  assign tmp2229 = (tmp2226 & tmp2227) | (tmp2226 & tmp2228) | (tmp2227 & tmp2228);
  wire tmp2230;
  assign tmp2230 = 1'b0;
  wire tmp2231;
  assign tmp2231 = 1'b0;
  wire tmp2232;
  assign tmp2232 = 1'b0;
  wire tmp2233;
  assign tmp2233 = (tmp2230 & tmp2231) | (tmp2230 & tmp2232) | (tmp2231 & tmp2232);
  wire tmp2234;
  assign tmp2234 = 1'b0;
  wire tmp2235;
  assign tmp2235 = 1'b0;
  wire tmp2236;
  assign tmp2236 = 1'b0;
  wire tmp2237;
  assign tmp2237 = (tmp2234 & tmp2235) | (tmp2234 & tmp2236) | (tmp2235 & tmp2236);
  wire tmp2238;
  assign tmp2238 = (tmp2229 & tmp2233) | (tmp2229 & tmp2237) | (tmp2233 & tmp2237);
  wire tmp2239;
  assign tmp2239 = 1'b0;
  wire tmp2240;
  assign tmp2240 = 1'b0;
  wire tmp2241;
  assign tmp2241 = 1'b0;
  wire tmp2242;
  assign tmp2242 = (tmp2239 & tmp2240) | (tmp2239 & tmp2241) | (tmp2240 & tmp2241);
  wire tmp2243;
  assign tmp2243 = 1'b0;
  wire tmp2244;
  assign tmp2244 = 1'b1;
  wire tmp2245;
  assign tmp2245 = 1'b0;
  wire tmp2246;
  assign tmp2246 = (tmp2243 & tmp2244) | (tmp2243 & tmp2245) | (tmp2244 & tmp2245);
  wire tmp2247;
  assign tmp2247 = 1'b0;
  wire tmp2248;
  assign tmp2248 = 1'b0;
  wire tmp2249;
  assign tmp2249 = 1'b0;
  wire tmp2250;
  assign tmp2250 = (tmp2247 & tmp2248) | (tmp2247 & tmp2249) | (tmp2248 & tmp2249);
  wire tmp2251;
  assign tmp2251 = (tmp2242 & tmp2246) | (tmp2242 & tmp2250) | (tmp2246 & tmp2250);
  wire tmp2252;
  assign tmp2252 = 1'b0;
  wire tmp2253;
  assign tmp2253 = 1'b0;
  wire tmp2254;
  assign tmp2254 = 1'b0;
  wire tmp2255;
  assign tmp2255 = (tmp2252 & tmp2253) | (tmp2252 & tmp2254) | (tmp2253 & tmp2254);
  wire tmp2256;
  assign tmp2256 = 1'b0;
  wire tmp2257;
  assign tmp2257 = 1'b0;
  wire tmp2258;
  assign tmp2258 = 1'b0;
  wire tmp2259;
  assign tmp2259 = (tmp2256 & tmp2257) | (tmp2256 & tmp2258) | (tmp2257 & tmp2258);
  wire tmp2260;
  assign tmp2260 = 1'b0;
  wire tmp2261;
  assign tmp2261 = 1'b0;
  wire tmp2262;
  assign tmp2262 = 1'b0;
  wire tmp2263;
  assign tmp2263 = (tmp2260 & tmp2261) | (tmp2260 & tmp2262) | (tmp2261 & tmp2262);
  wire tmp2264;
  assign tmp2264 = (tmp2255 & tmp2259) | (tmp2255 & tmp2263) | (tmp2259 & tmp2263);
  wire tmp2265;
  assign tmp2265 = (tmp2238 & tmp2251) | (tmp2238 & tmp2264) | (tmp2251 & tmp2264);
  wire tmp2266;
  assign tmp2266 = 1'b0;
  wire tmp2267;
  assign tmp2267 = 1'b0;
  wire tmp2268;
  assign tmp2268 = 1'b0;
  wire tmp2269;
  assign tmp2269 = (tmp2266 & tmp2267) | (tmp2266 & tmp2268) | (tmp2267 & tmp2268);
  wire tmp2270;
  assign tmp2270 = 1'b0;
  wire tmp2271;
  assign tmp2271 = 1'b0;
  wire tmp2272;
  assign tmp2272 = 1'b0;
  wire tmp2273;
  assign tmp2273 = (tmp2270 & tmp2271) | (tmp2270 & tmp2272) | (tmp2271 & tmp2272);
  wire tmp2274;
  assign tmp2274 = 1'b0;
  wire tmp2275;
  assign tmp2275 = 1'b0;
  wire tmp2276;
  assign tmp2276 = 1'b0;
  wire tmp2277;
  assign tmp2277 = (tmp2274 & tmp2275) | (tmp2274 & tmp2276) | (tmp2275 & tmp2276);
  wire tmp2278;
  assign tmp2278 = (tmp2269 & tmp2273) | (tmp2269 & tmp2277) | (tmp2273 & tmp2277);
  wire tmp2279;
  assign tmp2279 = 1'b0;
  wire tmp2280;
  assign tmp2280 = 1'b0;
  wire tmp2281;
  assign tmp2281 = 1'b0;
  wire tmp2282;
  assign tmp2282 = (tmp2279 & tmp2280) | (tmp2279 & tmp2281) | (tmp2280 & tmp2281);
  wire tmp2283;
  assign tmp2283 = 1'b0;
  wire tmp2284;
  assign tmp2284 = 1'b0;
  wire tmp2285;
  assign tmp2285 = 1'b0;
  wire tmp2286;
  assign tmp2286 = (tmp2283 & tmp2284) | (tmp2283 & tmp2285) | (tmp2284 & tmp2285);
  wire tmp2287;
  assign tmp2287 = 1'b0;
  wire tmp2288;
  assign tmp2288 = 1'b0;
  wire tmp2289;
  assign tmp2289 = 1'b0;
  wire tmp2290;
  assign tmp2290 = (tmp2287 & tmp2288) | (tmp2287 & tmp2289) | (tmp2288 & tmp2289);
  wire tmp2291;
  assign tmp2291 = (tmp2282 & tmp2286) | (tmp2282 & tmp2290) | (tmp2286 & tmp2290);
  wire tmp2292;
  assign tmp2292 = 1'b0;
  wire tmp2293;
  assign tmp2293 = 1'b0;
  wire tmp2294;
  assign tmp2294 = 1'b0;
  wire tmp2295;
  assign tmp2295 = (tmp2292 & tmp2293) | (tmp2292 & tmp2294) | (tmp2293 & tmp2294);
  wire tmp2296;
  assign tmp2296 = 1'b0;
  wire tmp2297;
  assign tmp2297 = 1'b0;
  wire tmp2298;
  assign tmp2298 = 1'b0;
  wire tmp2299;
  assign tmp2299 = (tmp2296 & tmp2297) | (tmp2296 & tmp2298) | (tmp2297 & tmp2298);
  wire tmp2300;
  assign tmp2300 = 1'b0;
  wire tmp2301;
  assign tmp2301 = 1'b0;
  wire tmp2302;
  assign tmp2302 = 1'b0;
  wire tmp2303;
  assign tmp2303 = (tmp2300 & tmp2301) | (tmp2300 & tmp2302) | (tmp2301 & tmp2302);
  wire tmp2304;
  assign tmp2304 = (tmp2295 & tmp2299) | (tmp2295 & tmp2303) | (tmp2299 & tmp2303);
  wire tmp2305;
  assign tmp2305 = (tmp2278 & tmp2291) | (tmp2278 & tmp2304) | (tmp2291 & tmp2304);
  wire tmp2306;
  assign tmp2306 = (tmp2225 & tmp2265) | (tmp2225 & tmp2305) | (tmp2265 & tmp2305);
  wire tmp2307;
  assign tmp2307 = 1'b0;
  wire tmp2308;
  assign tmp2308 = 1'b0;
  wire tmp2309;
  assign tmp2309 = 1'b0;
  wire tmp2310;
  assign tmp2310 = (tmp2307 & tmp2308) | (tmp2307 & tmp2309) | (tmp2308 & tmp2309);
  wire tmp2311;
  assign tmp2311 = 1'b0;
  wire tmp2312;
  assign tmp2312 = 1'b0;
  wire tmp2313;
  assign tmp2313 = 1'b0;
  wire tmp2314;
  assign tmp2314 = (tmp2311 & tmp2312) | (tmp2311 & tmp2313) | (tmp2312 & tmp2313);
  wire tmp2315;
  assign tmp2315 = 1'b0;
  wire tmp2316;
  assign tmp2316 = 1'b0;
  wire tmp2317;
  assign tmp2317 = 1'b0;
  wire tmp2318;
  assign tmp2318 = (tmp2315 & tmp2316) | (tmp2315 & tmp2317) | (tmp2316 & tmp2317);
  wire tmp2319;
  assign tmp2319 = (tmp2310 & tmp2314) | (tmp2310 & tmp2318) | (tmp2314 & tmp2318);
  wire tmp2320;
  assign tmp2320 = 1'b0;
  wire tmp2321;
  assign tmp2321 = 1'b0;
  wire tmp2322;
  assign tmp2322 = 1'b0;
  wire tmp2323;
  assign tmp2323 = (tmp2320 & tmp2321) | (tmp2320 & tmp2322) | (tmp2321 & tmp2322);
  wire tmp2324;
  assign tmp2324 = 1'b0;
  wire tmp2325;
  assign tmp2325 = 1'b1;
  wire tmp2326;
  assign tmp2326 = 1'b0;
  wire tmp2327;
  assign tmp2327 = (tmp2324 & tmp2325) | (tmp2324 & tmp2326) | (tmp2325 & tmp2326);
  wire tmp2328;
  assign tmp2328 = 1'b0;
  wire tmp2329;
  assign tmp2329 = 1'b0;
  wire tmp2330;
  assign tmp2330 = 1'b0;
  wire tmp2331;
  assign tmp2331 = (tmp2328 & tmp2329) | (tmp2328 & tmp2330) | (tmp2329 & tmp2330);
  wire tmp2332;
  assign tmp2332 = (tmp2323 & tmp2327) | (tmp2323 & tmp2331) | (tmp2327 & tmp2331);
  wire tmp2333;
  assign tmp2333 = 1'b0;
  wire tmp2334;
  assign tmp2334 = 1'b0;
  wire tmp2335;
  assign tmp2335 = 1'b0;
  wire tmp2336;
  assign tmp2336 = (tmp2333 & tmp2334) | (tmp2333 & tmp2335) | (tmp2334 & tmp2335);
  wire tmp2337;
  assign tmp2337 = 1'b0;
  wire tmp2338;
  assign tmp2338 = 1'b0;
  wire tmp2339;
  assign tmp2339 = 1'b0;
  wire tmp2340;
  assign tmp2340 = (tmp2337 & tmp2338) | (tmp2337 & tmp2339) | (tmp2338 & tmp2339);
  wire tmp2341;
  assign tmp2341 = 1'b0;
  wire tmp2342;
  assign tmp2342 = 1'b0;
  wire tmp2343;
  assign tmp2343 = 1'b0;
  wire tmp2344;
  assign tmp2344 = (tmp2341 & tmp2342) | (tmp2341 & tmp2343) | (tmp2342 & tmp2343);
  wire tmp2345;
  assign tmp2345 = (tmp2336 & tmp2340) | (tmp2336 & tmp2344) | (tmp2340 & tmp2344);
  wire tmp2346;
  assign tmp2346 = (tmp2319 & tmp2332) | (tmp2319 & tmp2345) | (tmp2332 & tmp2345);
  wire tmp2347;
  assign tmp2347 = 1'b0;
  wire tmp2348;
  assign tmp2348 = 1'b0;
  wire tmp2349;
  assign tmp2349 = 1'b0;
  wire tmp2350;
  assign tmp2350 = (tmp2347 & tmp2348) | (tmp2347 & tmp2349) | (tmp2348 & tmp2349);
  wire tmp2351;
  assign tmp2351 = 1'b0;
  wire tmp2352;
  assign tmp2352 = 1'b1;
  wire tmp2353;
  assign tmp2353 = 1'b0;
  wire tmp2354;
  assign tmp2354 = (tmp2351 & tmp2352) | (tmp2351 & tmp2353) | (tmp2352 & tmp2353);
  wire tmp2355;
  assign tmp2355 = 1'b0;
  wire tmp2356;
  assign tmp2356 = 1'b0;
  wire tmp2357;
  assign tmp2357 = 1'b0;
  wire tmp2358;
  assign tmp2358 = (tmp2355 & tmp2356) | (tmp2355 & tmp2357) | (tmp2356 & tmp2357);
  wire tmp2359;
  assign tmp2359 = (tmp2350 & tmp2354) | (tmp2350 & tmp2358) | (tmp2354 & tmp2358);
  wire tmp2360;
  assign tmp2360 = 1'b0;
  wire tmp2361;
  assign tmp2361 = 1'b1;
  wire tmp2362;
  assign tmp2362 = 1'b0;
  wire tmp2363;
  assign tmp2363 = (tmp2360 & tmp2361) | (tmp2360 & tmp2362) | (tmp2361 & tmp2362);
  wire tmp2364;
  assign tmp2364 = 1'b1;
  wire tmp2365;
  assign tmp2365 = 1'b1;
  wire tmp2366;
  assign tmp2366 = 1'b1;
  wire tmp2367;
  assign tmp2367 = (tmp2364 & tmp2365) | (tmp2364 & tmp2366) | (tmp2365 & tmp2366);
  wire tmp2368;
  assign tmp2368 = 1'b0;
  wire tmp2369;
  assign tmp2369 = 1'b1;
  wire tmp2370;
  assign tmp2370 = 1'b0;
  wire tmp2371;
  assign tmp2371 = (tmp2368 & tmp2369) | (tmp2368 & tmp2370) | (tmp2369 & tmp2370);
  wire tmp2372;
  assign tmp2372 = (tmp2363 & tmp2367) | (tmp2363 & tmp2371) | (tmp2367 & tmp2371);
  wire tmp2373;
  assign tmp2373 = 1'b0;
  wire tmp2374;
  assign tmp2374 = 1'b0;
  wire tmp2375;
  assign tmp2375 = 1'b0;
  wire tmp2376;
  assign tmp2376 = (tmp2373 & tmp2374) | (tmp2373 & tmp2375) | (tmp2374 & tmp2375);
  wire tmp2377;
  assign tmp2377 = 1'b0;
  wire tmp2378;
  assign tmp2378 = 1'b1;
  wire tmp2379;
  assign tmp2379 = 1'b0;
  wire tmp2380;
  assign tmp2380 = (tmp2377 & tmp2378) | (tmp2377 & tmp2379) | (tmp2378 & tmp2379);
  wire tmp2381;
  assign tmp2381 = 1'b0;
  wire tmp2382;
  assign tmp2382 = 1'b0;
  wire tmp2383;
  assign tmp2383 = 1'b0;
  wire tmp2384;
  assign tmp2384 = (tmp2381 & tmp2382) | (tmp2381 & tmp2383) | (tmp2382 & tmp2383);
  wire tmp2385;
  assign tmp2385 = (tmp2376 & tmp2380) | (tmp2376 & tmp2384) | (tmp2380 & tmp2384);
  wire tmp2386;
  assign tmp2386 = (tmp2359 & tmp2372) | (tmp2359 & tmp2385) | (tmp2372 & tmp2385);
  wire tmp2387;
  assign tmp2387 = 1'b0;
  wire tmp2388;
  assign tmp2388 = 1'b0;
  wire tmp2389;
  assign tmp2389 = 1'b0;
  wire tmp2390;
  assign tmp2390 = (tmp2387 & tmp2388) | (tmp2387 & tmp2389) | (tmp2388 & tmp2389);
  wire tmp2391;
  assign tmp2391 = 1'b0;
  wire tmp2392;
  assign tmp2392 = 1'b0;
  wire tmp2393;
  assign tmp2393 = 1'b0;
  wire tmp2394;
  assign tmp2394 = (tmp2391 & tmp2392) | (tmp2391 & tmp2393) | (tmp2392 & tmp2393);
  wire tmp2395;
  assign tmp2395 = 1'b0;
  wire tmp2396;
  assign tmp2396 = 1'b0;
  wire tmp2397;
  assign tmp2397 = 1'b0;
  wire tmp2398;
  assign tmp2398 = (tmp2395 & tmp2396) | (tmp2395 & tmp2397) | (tmp2396 & tmp2397);
  wire tmp2399;
  assign tmp2399 = (tmp2390 & tmp2394) | (tmp2390 & tmp2398) | (tmp2394 & tmp2398);
  wire tmp2400;
  assign tmp2400 = 1'b0;
  wire tmp2401;
  assign tmp2401 = 1'b0;
  wire tmp2402;
  assign tmp2402 = 1'b0;
  wire tmp2403;
  assign tmp2403 = (tmp2400 & tmp2401) | (tmp2400 & tmp2402) | (tmp2401 & tmp2402);
  wire tmp2404;
  assign tmp2404 = 1'b0;
  wire tmp2405;
  assign tmp2405 = 1'b1;
  wire tmp2406;
  assign tmp2406 = 1'b0;
  wire tmp2407;
  assign tmp2407 = (tmp2404 & tmp2405) | (tmp2404 & tmp2406) | (tmp2405 & tmp2406);
  wire tmp2408;
  assign tmp2408 = 1'b0;
  wire tmp2409;
  assign tmp2409 = 1'b0;
  wire tmp2410;
  assign tmp2410 = 1'b0;
  wire tmp2411;
  assign tmp2411 = (tmp2408 & tmp2409) | (tmp2408 & tmp2410) | (tmp2409 & tmp2410);
  wire tmp2412;
  assign tmp2412 = (tmp2403 & tmp2407) | (tmp2403 & tmp2411) | (tmp2407 & tmp2411);
  wire tmp2413;
  assign tmp2413 = 1'b0;
  wire tmp2414;
  assign tmp2414 = 1'b0;
  wire tmp2415;
  assign tmp2415 = 1'b0;
  wire tmp2416;
  assign tmp2416 = (tmp2413 & tmp2414) | (tmp2413 & tmp2415) | (tmp2414 & tmp2415);
  wire tmp2417;
  assign tmp2417 = 1'b0;
  wire tmp2418;
  assign tmp2418 = 1'b0;
  wire tmp2419;
  assign tmp2419 = 1'b0;
  wire tmp2420;
  assign tmp2420 = (tmp2417 & tmp2418) | (tmp2417 & tmp2419) | (tmp2418 & tmp2419);
  wire tmp2421;
  assign tmp2421 = 1'b0;
  wire tmp2422;
  assign tmp2422 = 1'b0;
  wire tmp2423;
  assign tmp2423 = 1'b0;
  wire tmp2424;
  assign tmp2424 = (tmp2421 & tmp2422) | (tmp2421 & tmp2423) | (tmp2422 & tmp2423);
  wire tmp2425;
  assign tmp2425 = (tmp2416 & tmp2420) | (tmp2416 & tmp2424) | (tmp2420 & tmp2424);
  wire tmp2426;
  assign tmp2426 = (tmp2399 & tmp2412) | (tmp2399 & tmp2425) | (tmp2412 & tmp2425);
  wire tmp2427;
  assign tmp2427 = (tmp2346 & tmp2386) | (tmp2346 & tmp2426) | (tmp2386 & tmp2426);
  wire tmp2428;
  assign tmp2428 = 1'b0;
  wire tmp2429;
  assign tmp2429 = 1'b0;
  wire tmp2430;
  assign tmp2430 = 1'b0;
  wire tmp2431;
  assign tmp2431 = (tmp2428 & tmp2429) | (tmp2428 & tmp2430) | (tmp2429 & tmp2430);
  wire tmp2432;
  assign tmp2432 = 1'b0;
  wire tmp2433;
  assign tmp2433 = 1'b0;
  wire tmp2434;
  assign tmp2434 = 1'b0;
  wire tmp2435;
  assign tmp2435 = (tmp2432 & tmp2433) | (tmp2432 & tmp2434) | (tmp2433 & tmp2434);
  wire tmp2436;
  assign tmp2436 = 1'b0;
  wire tmp2437;
  assign tmp2437 = 1'b0;
  wire tmp2438;
  assign tmp2438 = 1'b0;
  wire tmp2439;
  assign tmp2439 = (tmp2436 & tmp2437) | (tmp2436 & tmp2438) | (tmp2437 & tmp2438);
  wire tmp2440;
  assign tmp2440 = (tmp2431 & tmp2435) | (tmp2431 & tmp2439) | (tmp2435 & tmp2439);
  wire tmp2441;
  assign tmp2441 = 1'b0;
  wire tmp2442;
  assign tmp2442 = 1'b0;
  wire tmp2443;
  assign tmp2443 = 1'b0;
  wire tmp2444;
  assign tmp2444 = (tmp2441 & tmp2442) | (tmp2441 & tmp2443) | (tmp2442 & tmp2443);
  wire tmp2445;
  assign tmp2445 = 1'b0;
  wire tmp2446;
  assign tmp2446 = 1'b0;
  wire tmp2447;
  assign tmp2447 = 1'b0;
  wire tmp2448;
  assign tmp2448 = (tmp2445 & tmp2446) | (tmp2445 & tmp2447) | (tmp2446 & tmp2447);
  wire tmp2449;
  assign tmp2449 = 1'b0;
  wire tmp2450;
  assign tmp2450 = 1'b0;
  wire tmp2451;
  assign tmp2451 = 1'b0;
  wire tmp2452;
  assign tmp2452 = (tmp2449 & tmp2450) | (tmp2449 & tmp2451) | (tmp2450 & tmp2451);
  wire tmp2453;
  assign tmp2453 = (tmp2444 & tmp2448) | (tmp2444 & tmp2452) | (tmp2448 & tmp2452);
  wire tmp2454;
  assign tmp2454 = 1'b0;
  wire tmp2455;
  assign tmp2455 = 1'b0;
  wire tmp2456;
  assign tmp2456 = 1'b0;
  wire tmp2457;
  assign tmp2457 = (tmp2454 & tmp2455) | (tmp2454 & tmp2456) | (tmp2455 & tmp2456);
  wire tmp2458;
  assign tmp2458 = 1'b0;
  wire tmp2459;
  assign tmp2459 = 1'b0;
  wire tmp2460;
  assign tmp2460 = 1'b0;
  wire tmp2461;
  assign tmp2461 = (tmp2458 & tmp2459) | (tmp2458 & tmp2460) | (tmp2459 & tmp2460);
  wire tmp2462;
  assign tmp2462 = 1'b0;
  wire tmp2463;
  assign tmp2463 = 1'b0;
  wire tmp2464;
  assign tmp2464 = 1'b0;
  wire tmp2465;
  assign tmp2465 = (tmp2462 & tmp2463) | (tmp2462 & tmp2464) | (tmp2463 & tmp2464);
  wire tmp2466;
  assign tmp2466 = (tmp2457 & tmp2461) | (tmp2457 & tmp2465) | (tmp2461 & tmp2465);
  wire tmp2467;
  assign tmp2467 = (tmp2440 & tmp2453) | (tmp2440 & tmp2466) | (tmp2453 & tmp2466);
  wire tmp2468;
  assign tmp2468 = 1'b0;
  wire tmp2469;
  assign tmp2469 = 1'b0;
  wire tmp2470;
  assign tmp2470 = 1'b0;
  wire tmp2471;
  assign tmp2471 = (tmp2468 & tmp2469) | (tmp2468 & tmp2470) | (tmp2469 & tmp2470);
  wire tmp2472;
  assign tmp2472 = 1'b0;
  wire tmp2473;
  assign tmp2473 = 1'b0;
  wire tmp2474;
  assign tmp2474 = 1'b0;
  wire tmp2475;
  assign tmp2475 = (tmp2472 & tmp2473) | (tmp2472 & tmp2474) | (tmp2473 & tmp2474);
  wire tmp2476;
  assign tmp2476 = 1'b0;
  wire tmp2477;
  assign tmp2477 = 1'b0;
  wire tmp2478;
  assign tmp2478 = 1'b0;
  wire tmp2479;
  assign tmp2479 = (tmp2476 & tmp2477) | (tmp2476 & tmp2478) | (tmp2477 & tmp2478);
  wire tmp2480;
  assign tmp2480 = (tmp2471 & tmp2475) | (tmp2471 & tmp2479) | (tmp2475 & tmp2479);
  wire tmp2481;
  assign tmp2481 = 1'b0;
  wire tmp2482;
  assign tmp2482 = 1'b0;
  wire tmp2483;
  assign tmp2483 = 1'b0;
  wire tmp2484;
  assign tmp2484 = (tmp2481 & tmp2482) | (tmp2481 & tmp2483) | (tmp2482 & tmp2483);
  wire tmp2485;
  assign tmp2485 = 1'b0;
  wire tmp2486;
  assign tmp2486 = 1'b1;
  wire tmp2487;
  assign tmp2487 = 1'b0;
  wire tmp2488;
  assign tmp2488 = (tmp2485 & tmp2486) | (tmp2485 & tmp2487) | (tmp2486 & tmp2487);
  wire tmp2489;
  assign tmp2489 = 1'b0;
  wire tmp2490;
  assign tmp2490 = 1'b0;
  wire tmp2491;
  assign tmp2491 = 1'b0;
  wire tmp2492;
  assign tmp2492 = (tmp2489 & tmp2490) | (tmp2489 & tmp2491) | (tmp2490 & tmp2491);
  wire tmp2493;
  assign tmp2493 = (tmp2484 & tmp2488) | (tmp2484 & tmp2492) | (tmp2488 & tmp2492);
  wire tmp2494;
  assign tmp2494 = 1'b0;
  wire tmp2495;
  assign tmp2495 = 1'b0;
  wire tmp2496;
  assign tmp2496 = 1'b0;
  wire tmp2497;
  assign tmp2497 = (tmp2494 & tmp2495) | (tmp2494 & tmp2496) | (tmp2495 & tmp2496);
  wire tmp2498;
  assign tmp2498 = 1'b0;
  wire tmp2499;
  assign tmp2499 = 1'b0;
  wire tmp2500;
  assign tmp2500 = 1'b0;
  wire tmp2501;
  assign tmp2501 = (tmp2498 & tmp2499) | (tmp2498 & tmp2500) | (tmp2499 & tmp2500);
  wire tmp2502;
  assign tmp2502 = 1'b0;
  wire tmp2503;
  assign tmp2503 = 1'b0;
  wire tmp2504;
  assign tmp2504 = 1'b0;
  wire tmp2505;
  assign tmp2505 = (tmp2502 & tmp2503) | (tmp2502 & tmp2504) | (tmp2503 & tmp2504);
  wire tmp2506;
  assign tmp2506 = (tmp2497 & tmp2501) | (tmp2497 & tmp2505) | (tmp2501 & tmp2505);
  wire tmp2507;
  assign tmp2507 = (tmp2480 & tmp2493) | (tmp2480 & tmp2506) | (tmp2493 & tmp2506);
  wire tmp2508;
  assign tmp2508 = 1'b0;
  wire tmp2509;
  assign tmp2509 = 1'b0;
  wire tmp2510;
  assign tmp2510 = 1'b0;
  wire tmp2511;
  assign tmp2511 = (tmp2508 & tmp2509) | (tmp2508 & tmp2510) | (tmp2509 & tmp2510);
  wire tmp2512;
  assign tmp2512 = 1'b0;
  wire tmp2513;
  assign tmp2513 = 1'b0;
  wire tmp2514;
  assign tmp2514 = 1'b0;
  wire tmp2515;
  assign tmp2515 = (tmp2512 & tmp2513) | (tmp2512 & tmp2514) | (tmp2513 & tmp2514);
  wire tmp2516;
  assign tmp2516 = 1'b0;
  wire tmp2517;
  assign tmp2517 = 1'b0;
  wire tmp2518;
  assign tmp2518 = 1'b0;
  wire tmp2519;
  assign tmp2519 = (tmp2516 & tmp2517) | (tmp2516 & tmp2518) | (tmp2517 & tmp2518);
  wire tmp2520;
  assign tmp2520 = (tmp2511 & tmp2515) | (tmp2511 & tmp2519) | (tmp2515 & tmp2519);
  wire tmp2521;
  assign tmp2521 = 1'b0;
  wire tmp2522;
  assign tmp2522 = 1'b0;
  wire tmp2523;
  assign tmp2523 = 1'b0;
  wire tmp2524;
  assign tmp2524 = (tmp2521 & tmp2522) | (tmp2521 & tmp2523) | (tmp2522 & tmp2523);
  wire tmp2525;
  assign tmp2525 = 1'b0;
  wire tmp2526;
  assign tmp2526 = 1'b0;
  wire tmp2527;
  assign tmp2527 = 1'b0;
  wire tmp2528;
  assign tmp2528 = (tmp2525 & tmp2526) | (tmp2525 & tmp2527) | (tmp2526 & tmp2527);
  wire tmp2529;
  assign tmp2529 = 1'b0;
  wire tmp2530;
  assign tmp2530 = 1'b0;
  wire tmp2531;
  assign tmp2531 = 1'b0;
  wire tmp2532;
  assign tmp2532 = (tmp2529 & tmp2530) | (tmp2529 & tmp2531) | (tmp2530 & tmp2531);
  wire tmp2533;
  assign tmp2533 = (tmp2524 & tmp2528) | (tmp2524 & tmp2532) | (tmp2528 & tmp2532);
  wire tmp2534;
  assign tmp2534 = 1'b0;
  wire tmp2535;
  assign tmp2535 = 1'b0;
  wire tmp2536;
  assign tmp2536 = 1'b0;
  wire tmp2537;
  assign tmp2537 = (tmp2534 & tmp2535) | (tmp2534 & tmp2536) | (tmp2535 & tmp2536);
  wire tmp2538;
  assign tmp2538 = 1'b0;
  wire tmp2539;
  assign tmp2539 = 1'b0;
  wire tmp2540;
  assign tmp2540 = 1'b0;
  wire tmp2541;
  assign tmp2541 = (tmp2538 & tmp2539) | (tmp2538 & tmp2540) | (tmp2539 & tmp2540);
  wire tmp2542;
  assign tmp2542 = 1'b0;
  wire tmp2543;
  assign tmp2543 = 1'b0;
  wire tmp2544;
  assign tmp2544 = 1'b0;
  wire tmp2545;
  assign tmp2545 = (tmp2542 & tmp2543) | (tmp2542 & tmp2544) | (tmp2543 & tmp2544);
  wire tmp2546;
  assign tmp2546 = (tmp2537 & tmp2541) | (tmp2537 & tmp2545) | (tmp2541 & tmp2545);
  wire tmp2547;
  assign tmp2547 = (tmp2520 & tmp2533) | (tmp2520 & tmp2546) | (tmp2533 & tmp2546);
  wire tmp2548;
  assign tmp2548 = (tmp2467 & tmp2507) | (tmp2467 & tmp2547) | (tmp2507 & tmp2547);
  wire tmp2549;
  assign tmp2549 = (tmp2306 & tmp2427) | (tmp2306 & tmp2548) | (tmp2427 & tmp2548);
  wire tmp2550;
  assign tmp2550 = 1'b0;
  wire tmp2551;
  assign tmp2551 = 1'b0;
  wire tmp2552;
  assign tmp2552 = 1'b0;
  wire tmp2553;
  assign tmp2553 = (tmp2550 & tmp2551) | (tmp2550 & tmp2552) | (tmp2551 & tmp2552);
  wire tmp2554;
  assign tmp2554 = 1'b0;
  wire tmp2555;
  assign tmp2555 = 1'b0;
  wire tmp2556;
  assign tmp2556 = 1'b0;
  wire tmp2557;
  assign tmp2557 = (tmp2554 & tmp2555) | (tmp2554 & tmp2556) | (tmp2555 & tmp2556);
  wire tmp2558;
  assign tmp2558 = 1'b0;
  wire tmp2559;
  assign tmp2559 = 1'b0;
  wire tmp2560;
  assign tmp2560 = 1'b0;
  wire tmp2561;
  assign tmp2561 = (tmp2558 & tmp2559) | (tmp2558 & tmp2560) | (tmp2559 & tmp2560);
  wire tmp2562;
  assign tmp2562 = (tmp2553 & tmp2557) | (tmp2553 & tmp2561) | (tmp2557 & tmp2561);
  wire tmp2563;
  assign tmp2563 = 1'b0;
  wire tmp2564;
  assign tmp2564 = 1'b0;
  wire tmp2565;
  assign tmp2565 = 1'b0;
  wire tmp2566;
  assign tmp2566 = (tmp2563 & tmp2564) | (tmp2563 & tmp2565) | (tmp2564 & tmp2565);
  wire tmp2567;
  assign tmp2567 = 1'b0;
  wire tmp2568;
  assign tmp2568 = 1'b1;
  wire tmp2569;
  assign tmp2569 = 1'b0;
  wire tmp2570;
  assign tmp2570 = (tmp2567 & tmp2568) | (tmp2567 & tmp2569) | (tmp2568 & tmp2569);
  wire tmp2571;
  assign tmp2571 = 1'b0;
  wire tmp2572;
  assign tmp2572 = 1'b0;
  wire tmp2573;
  assign tmp2573 = 1'b0;
  wire tmp2574;
  assign tmp2574 = (tmp2571 & tmp2572) | (tmp2571 & tmp2573) | (tmp2572 & tmp2573);
  wire tmp2575;
  assign tmp2575 = (tmp2566 & tmp2570) | (tmp2566 & tmp2574) | (tmp2570 & tmp2574);
  wire tmp2576;
  assign tmp2576 = 1'b0;
  wire tmp2577;
  assign tmp2577 = 1'b0;
  wire tmp2578;
  assign tmp2578 = 1'b0;
  wire tmp2579;
  assign tmp2579 = (tmp2576 & tmp2577) | (tmp2576 & tmp2578) | (tmp2577 & tmp2578);
  wire tmp2580;
  assign tmp2580 = 1'b0;
  wire tmp2581;
  assign tmp2581 = 1'b0;
  wire tmp2582;
  assign tmp2582 = 1'b0;
  wire tmp2583;
  assign tmp2583 = (tmp2580 & tmp2581) | (tmp2580 & tmp2582) | (tmp2581 & tmp2582);
  wire tmp2584;
  assign tmp2584 = 1'b0;
  wire tmp2585;
  assign tmp2585 = 1'b0;
  wire tmp2586;
  assign tmp2586 = 1'b0;
  wire tmp2587;
  assign tmp2587 = (tmp2584 & tmp2585) | (tmp2584 & tmp2586) | (tmp2585 & tmp2586);
  wire tmp2588;
  assign tmp2588 = (tmp2579 & tmp2583) | (tmp2579 & tmp2587) | (tmp2583 & tmp2587);
  wire tmp2589;
  assign tmp2589 = (tmp2562 & tmp2575) | (tmp2562 & tmp2588) | (tmp2575 & tmp2588);
  wire tmp2590;
  assign tmp2590 = 1'b0;
  wire tmp2591;
  assign tmp2591 = 1'b0;
  wire tmp2592;
  assign tmp2592 = 1'b0;
  wire tmp2593;
  assign tmp2593 = (tmp2590 & tmp2591) | (tmp2590 & tmp2592) | (tmp2591 & tmp2592);
  wire tmp2594;
  assign tmp2594 = 1'b0;
  wire tmp2595;
  assign tmp2595 = 1'b1;
  wire tmp2596;
  assign tmp2596 = 1'b0;
  wire tmp2597;
  assign tmp2597 = (tmp2594 & tmp2595) | (tmp2594 & tmp2596) | (tmp2595 & tmp2596);
  wire tmp2598;
  assign tmp2598 = 1'b0;
  wire tmp2599;
  assign tmp2599 = 1'b0;
  wire tmp2600;
  assign tmp2600 = 1'b0;
  wire tmp2601;
  assign tmp2601 = (tmp2598 & tmp2599) | (tmp2598 & tmp2600) | (tmp2599 & tmp2600);
  wire tmp2602;
  assign tmp2602 = (tmp2593 & tmp2597) | (tmp2593 & tmp2601) | (tmp2597 & tmp2601);
  wire tmp2603;
  assign tmp2603 = 1'b0;
  wire tmp2604;
  assign tmp2604 = 1'b1;
  wire tmp2605;
  assign tmp2605 = 1'b0;
  wire tmp2606;
  assign tmp2606 = (tmp2603 & tmp2604) | (tmp2603 & tmp2605) | (tmp2604 & tmp2605);
  wire tmp2607;
  assign tmp2607 = 1'b1;
  wire tmp2608;
  assign tmp2608 = 1'b1;
  wire tmp2609;
  assign tmp2609 = 1'b1;
  wire tmp2610;
  assign tmp2610 = (tmp2607 & tmp2608) | (tmp2607 & tmp2609) | (tmp2608 & tmp2609);
  wire tmp2611;
  assign tmp2611 = 1'b0;
  wire tmp2612;
  assign tmp2612 = 1'b1;
  wire tmp2613;
  assign tmp2613 = 1'b0;
  wire tmp2614;
  assign tmp2614 = (tmp2611 & tmp2612) | (tmp2611 & tmp2613) | (tmp2612 & tmp2613);
  wire tmp2615;
  assign tmp2615 = (tmp2606 & tmp2610) | (tmp2606 & tmp2614) | (tmp2610 & tmp2614);
  wire tmp2616;
  assign tmp2616 = 1'b0;
  wire tmp2617;
  assign tmp2617 = 1'b0;
  wire tmp2618;
  assign tmp2618 = 1'b0;
  wire tmp2619;
  assign tmp2619 = (tmp2616 & tmp2617) | (tmp2616 & tmp2618) | (tmp2617 & tmp2618);
  wire tmp2620;
  assign tmp2620 = 1'b0;
  wire tmp2621;
  assign tmp2621 = 1'b1;
  wire tmp2622;
  assign tmp2622 = 1'b0;
  wire tmp2623;
  assign tmp2623 = (tmp2620 & tmp2621) | (tmp2620 & tmp2622) | (tmp2621 & tmp2622);
  wire tmp2624;
  assign tmp2624 = 1'b0;
  wire tmp2625;
  assign tmp2625 = 1'b0;
  wire tmp2626;
  assign tmp2626 = 1'b0;
  wire tmp2627;
  assign tmp2627 = (tmp2624 & tmp2625) | (tmp2624 & tmp2626) | (tmp2625 & tmp2626);
  wire tmp2628;
  assign tmp2628 = (tmp2619 & tmp2623) | (tmp2619 & tmp2627) | (tmp2623 & tmp2627);
  wire tmp2629;
  assign tmp2629 = (tmp2602 & tmp2615) | (tmp2602 & tmp2628) | (tmp2615 & tmp2628);
  wire tmp2630;
  assign tmp2630 = 1'b0;
  wire tmp2631;
  assign tmp2631 = 1'b0;
  wire tmp2632;
  assign tmp2632 = 1'b0;
  wire tmp2633;
  assign tmp2633 = (tmp2630 & tmp2631) | (tmp2630 & tmp2632) | (tmp2631 & tmp2632);
  wire tmp2634;
  assign tmp2634 = 1'b0;
  wire tmp2635;
  assign tmp2635 = 1'b0;
  wire tmp2636;
  assign tmp2636 = 1'b0;
  wire tmp2637;
  assign tmp2637 = (tmp2634 & tmp2635) | (tmp2634 & tmp2636) | (tmp2635 & tmp2636);
  wire tmp2638;
  assign tmp2638 = 1'b0;
  wire tmp2639;
  assign tmp2639 = 1'b0;
  wire tmp2640;
  assign tmp2640 = 1'b0;
  wire tmp2641;
  assign tmp2641 = (tmp2638 & tmp2639) | (tmp2638 & tmp2640) | (tmp2639 & tmp2640);
  wire tmp2642;
  assign tmp2642 = (tmp2633 & tmp2637) | (tmp2633 & tmp2641) | (tmp2637 & tmp2641);
  wire tmp2643;
  assign tmp2643 = 1'b0;
  wire tmp2644;
  assign tmp2644 = 1'b0;
  wire tmp2645;
  assign tmp2645 = 1'b0;
  wire tmp2646;
  assign tmp2646 = (tmp2643 & tmp2644) | (tmp2643 & tmp2645) | (tmp2644 & tmp2645);
  wire tmp2647;
  assign tmp2647 = 1'b0;
  wire tmp2648;
  assign tmp2648 = 1'b1;
  wire tmp2649;
  assign tmp2649 = 1'b0;
  wire tmp2650;
  assign tmp2650 = (tmp2647 & tmp2648) | (tmp2647 & tmp2649) | (tmp2648 & tmp2649);
  wire tmp2651;
  assign tmp2651 = 1'b0;
  wire tmp2652;
  assign tmp2652 = 1'b0;
  wire tmp2653;
  assign tmp2653 = 1'b0;
  wire tmp2654;
  assign tmp2654 = (tmp2651 & tmp2652) | (tmp2651 & tmp2653) | (tmp2652 & tmp2653);
  wire tmp2655;
  assign tmp2655 = (tmp2646 & tmp2650) | (tmp2646 & tmp2654) | (tmp2650 & tmp2654);
  wire tmp2656;
  assign tmp2656 = 1'b0;
  wire tmp2657;
  assign tmp2657 = 1'b0;
  wire tmp2658;
  assign tmp2658 = 1'b0;
  wire tmp2659;
  assign tmp2659 = (tmp2656 & tmp2657) | (tmp2656 & tmp2658) | (tmp2657 & tmp2658);
  wire tmp2660;
  assign tmp2660 = 1'b0;
  wire tmp2661;
  assign tmp2661 = 1'b0;
  wire tmp2662;
  assign tmp2662 = 1'b0;
  wire tmp2663;
  assign tmp2663 = (tmp2660 & tmp2661) | (tmp2660 & tmp2662) | (tmp2661 & tmp2662);
  wire tmp2664;
  assign tmp2664 = 1'b0;
  wire tmp2665;
  assign tmp2665 = 1'b0;
  wire tmp2666;
  assign tmp2666 = 1'b0;
  wire tmp2667;
  assign tmp2667 = (tmp2664 & tmp2665) | (tmp2664 & tmp2666) | (tmp2665 & tmp2666);
  wire tmp2668;
  assign tmp2668 = (tmp2659 & tmp2663) | (tmp2659 & tmp2667) | (tmp2663 & tmp2667);
  wire tmp2669;
  assign tmp2669 = (tmp2642 & tmp2655) | (tmp2642 & tmp2668) | (tmp2655 & tmp2668);
  wire tmp2670;
  assign tmp2670 = (tmp2589 & tmp2629) | (tmp2589 & tmp2669) | (tmp2629 & tmp2669);
  wire tmp2671;
  assign tmp2671 = 1'b0;
  wire tmp2672;
  assign tmp2672 = 1'b0;
  wire tmp2673;
  assign tmp2673 = 1'b0;
  wire tmp2674;
  assign tmp2674 = (tmp2671 & tmp2672) | (tmp2671 & tmp2673) | (tmp2672 & tmp2673);
  wire tmp2675;
  assign tmp2675 = 1'b0;
  wire tmp2676;
  assign tmp2676 = 1'b1;
  wire tmp2677;
  assign tmp2677 = 1'b0;
  wire tmp2678;
  assign tmp2678 = (tmp2675 & tmp2676) | (tmp2675 & tmp2677) | (tmp2676 & tmp2677);
  wire tmp2679;
  assign tmp2679 = 1'b0;
  wire tmp2680;
  assign tmp2680 = 1'b0;
  wire tmp2681;
  assign tmp2681 = 1'b0;
  wire tmp2682;
  assign tmp2682 = (tmp2679 & tmp2680) | (tmp2679 & tmp2681) | (tmp2680 & tmp2681);
  wire tmp2683;
  assign tmp2683 = (tmp2674 & tmp2678) | (tmp2674 & tmp2682) | (tmp2678 & tmp2682);
  wire tmp2684;
  assign tmp2684 = 1'b0;
  wire tmp2685;
  assign tmp2685 = 1'b1;
  wire tmp2686;
  assign tmp2686 = 1'b0;
  wire tmp2687;
  assign tmp2687 = (tmp2684 & tmp2685) | (tmp2684 & tmp2686) | (tmp2685 & tmp2686);
  wire tmp2688;
  assign tmp2688 = 1'b1;
  wire tmp2689;
  assign tmp2689 = 1'b1;
  wire tmp2690;
  assign tmp2690 = 1'b1;
  wire tmp2691;
  assign tmp2691 = (tmp2688 & tmp2689) | (tmp2688 & tmp2690) | (tmp2689 & tmp2690);
  wire tmp2692;
  assign tmp2692 = 1'b0;
  wire tmp2693;
  assign tmp2693 = 1'b1;
  wire tmp2694;
  assign tmp2694 = 1'b0;
  wire tmp2695;
  assign tmp2695 = (tmp2692 & tmp2693) | (tmp2692 & tmp2694) | (tmp2693 & tmp2694);
  wire tmp2696;
  assign tmp2696 = (tmp2687 & tmp2691) | (tmp2687 & tmp2695) | (tmp2691 & tmp2695);
  wire tmp2697;
  assign tmp2697 = 1'b0;
  wire tmp2698;
  assign tmp2698 = 1'b0;
  wire tmp2699;
  assign tmp2699 = 1'b0;
  wire tmp2700;
  assign tmp2700 = (tmp2697 & tmp2698) | (tmp2697 & tmp2699) | (tmp2698 & tmp2699);
  wire tmp2701;
  assign tmp2701 = 1'b0;
  wire tmp2702;
  assign tmp2702 = 1'b1;
  wire tmp2703;
  assign tmp2703 = 1'b0;
  wire tmp2704;
  assign tmp2704 = (tmp2701 & tmp2702) | (tmp2701 & tmp2703) | (tmp2702 & tmp2703);
  wire tmp2705;
  assign tmp2705 = 1'b0;
  wire tmp2706;
  assign tmp2706 = 1'b0;
  wire tmp2707;
  assign tmp2707 = 1'b0;
  wire tmp2708;
  assign tmp2708 = (tmp2705 & tmp2706) | (tmp2705 & tmp2707) | (tmp2706 & tmp2707);
  wire tmp2709;
  assign tmp2709 = (tmp2700 & tmp2704) | (tmp2700 & tmp2708) | (tmp2704 & tmp2708);
  wire tmp2710;
  assign tmp2710 = (tmp2683 & tmp2696) | (tmp2683 & tmp2709) | (tmp2696 & tmp2709);
  wire tmp2711;
  assign tmp2711 = 1'b0;
  wire tmp2712;
  assign tmp2712 = 1'b1;
  wire tmp2713;
  assign tmp2713 = 1'b0;
  wire tmp2714;
  assign tmp2714 = (tmp2711 & tmp2712) | (tmp2711 & tmp2713) | (tmp2712 & tmp2713);
  wire tmp2715;
  assign tmp2715 = 1'b1;
  wire tmp2716;
  assign tmp2716 = 1'b1;
  wire tmp2717;
  assign tmp2717 = 1'b1;
  wire tmp2718;
  assign tmp2718 = (tmp2715 & tmp2716) | (tmp2715 & tmp2717) | (tmp2716 & tmp2717);
  wire tmp2719;
  assign tmp2719 = 1'b0;
  wire tmp2720;
  assign tmp2720 = 1'b1;
  wire tmp2721;
  assign tmp2721 = 1'b0;
  wire tmp2722;
  assign tmp2722 = (tmp2719 & tmp2720) | (tmp2719 & tmp2721) | (tmp2720 & tmp2721);
  wire tmp2723;
  assign tmp2723 = (tmp2714 & tmp2718) | (tmp2714 & tmp2722) | (tmp2718 & tmp2722);
  wire tmp2724;
  assign tmp2724 = 1'b1;
  wire tmp2725;
  assign tmp2725 = 1'b1;
  wire tmp2726;
  assign tmp2726 = 1'b1;
  wire tmp2727;
  assign tmp2727 = (tmp2724 & tmp2725) | (tmp2724 & tmp2726) | (tmp2725 & tmp2726);
  wire tmp2728;
  assign tmp2728 = 1'b1;
  wire tmp2729;
  assign tmp2729 = ~pi5;
  wire tmp2730;
  assign tmp2730 = ~pi6;
  wire tmp2731;
  assign tmp2731 = (tmp2728 & tmp2729) | (tmp2728 & tmp2730) | (tmp2729 & tmp2730);
  wire tmp2732;
  assign tmp2732 = 1'b1;
  wire tmp2733;
  assign tmp2733 = ~pi6;
  wire tmp2734;
  assign tmp2734 = ~pi7;
  wire tmp2735;
  assign tmp2735 = (tmp2732 & tmp2733) | (tmp2732 & tmp2734) | (tmp2733 & tmp2734);
  wire tmp2736;
  assign tmp2736 = (tmp2727 & tmp2731) | (tmp2727 & tmp2735) | (tmp2731 & tmp2735);
  wire tmp2737;
  assign tmp2737 = 1'b0;
  wire tmp2738;
  assign tmp2738 = 1'b1;
  wire tmp2739;
  assign tmp2739 = 1'b0;
  wire tmp2740;
  assign tmp2740 = (tmp2737 & tmp2738) | (tmp2737 & tmp2739) | (tmp2738 & tmp2739);
  wire tmp2741;
  assign tmp2741 = 1'b1;
  wire tmp2742;
  assign tmp2742 = ~pi6;
  wire tmp2743;
  assign tmp2743 = ~pi7;
  wire tmp2744;
  assign tmp2744 = (tmp2741 & tmp2742) | (tmp2741 & tmp2743) | (tmp2742 & tmp2743);
  wire tmp2745;
  assign tmp2745 = 1'b0;
  wire tmp2746;
  assign tmp2746 = ~pi7;
  wire tmp2747;
  assign tmp2747 = 1'b0;
  wire tmp2748;
  assign tmp2748 = (tmp2745 & tmp2746) | (tmp2745 & tmp2747) | (tmp2746 & tmp2747);
  wire tmp2749;
  assign tmp2749 = (tmp2740 & tmp2744) | (tmp2740 & tmp2748) | (tmp2744 & tmp2748);
  wire tmp2750;
  assign tmp2750 = (tmp2723 & tmp2736) | (tmp2723 & tmp2749) | (tmp2736 & tmp2749);
  wire tmp2751;
  assign tmp2751 = 1'b0;
  wire tmp2752;
  assign tmp2752 = 1'b0;
  wire tmp2753;
  assign tmp2753 = 1'b0;
  wire tmp2754;
  assign tmp2754 = (tmp2751 & tmp2752) | (tmp2751 & tmp2753) | (tmp2752 & tmp2753);
  wire tmp2755;
  assign tmp2755 = 1'b0;
  wire tmp2756;
  assign tmp2756 = 1'b1;
  wire tmp2757;
  assign tmp2757 = 1'b0;
  wire tmp2758;
  assign tmp2758 = (tmp2755 & tmp2756) | (tmp2755 & tmp2757) | (tmp2756 & tmp2757);
  wire tmp2759;
  assign tmp2759 = 1'b0;
  wire tmp2760;
  assign tmp2760 = 1'b0;
  wire tmp2761;
  assign tmp2761 = 1'b0;
  wire tmp2762;
  assign tmp2762 = (tmp2759 & tmp2760) | (tmp2759 & tmp2761) | (tmp2760 & tmp2761);
  wire tmp2763;
  assign tmp2763 = (tmp2754 & tmp2758) | (tmp2754 & tmp2762) | (tmp2758 & tmp2762);
  wire tmp2764;
  assign tmp2764 = 1'b0;
  wire tmp2765;
  assign tmp2765 = 1'b1;
  wire tmp2766;
  assign tmp2766 = 1'b0;
  wire tmp2767;
  assign tmp2767 = (tmp2764 & tmp2765) | (tmp2764 & tmp2766) | (tmp2765 & tmp2766);
  wire tmp2768;
  assign tmp2768 = 1'b1;
  wire tmp2769;
  assign tmp2769 = ~pi6;
  wire tmp2770;
  assign tmp2770 = ~pi7;
  wire tmp2771;
  assign tmp2771 = (tmp2768 & tmp2769) | (tmp2768 & tmp2770) | (tmp2769 & tmp2770);
  wire tmp2772;
  assign tmp2772 = 1'b0;
  wire tmp2773;
  assign tmp2773 = ~pi7;
  wire tmp2774;
  assign tmp2774 = 1'b0;
  wire tmp2775;
  assign tmp2775 = (tmp2772 & tmp2773) | (tmp2772 & tmp2774) | (tmp2773 & tmp2774);
  wire tmp2776;
  assign tmp2776 = (tmp2767 & tmp2771) | (tmp2767 & tmp2775) | (tmp2771 & tmp2775);
  wire tmp2777;
  assign tmp2777 = 1'b0;
  wire tmp2778;
  assign tmp2778 = 1'b0;
  wire tmp2779;
  assign tmp2779 = 1'b0;
  wire tmp2780;
  assign tmp2780 = (tmp2777 & tmp2778) | (tmp2777 & tmp2779) | (tmp2778 & tmp2779);
  wire tmp2781;
  assign tmp2781 = 1'b0;
  wire tmp2782;
  assign tmp2782 = ~pi7;
  wire tmp2783;
  assign tmp2783 = 1'b0;
  wire tmp2784;
  assign tmp2784 = (tmp2781 & tmp2782) | (tmp2781 & tmp2783) | (tmp2782 & tmp2783);
  wire tmp2785;
  assign tmp2785 = 1'b0;
  wire tmp2786;
  assign tmp2786 = 1'b0;
  wire tmp2787;
  assign tmp2787 = 1'b0;
  wire tmp2788;
  assign tmp2788 = (tmp2785 & tmp2786) | (tmp2785 & tmp2787) | (tmp2786 & tmp2787);
  wire tmp2789;
  assign tmp2789 = (tmp2780 & tmp2784) | (tmp2780 & tmp2788) | (tmp2784 & tmp2788);
  wire tmp2790;
  assign tmp2790 = (tmp2763 & tmp2776) | (tmp2763 & tmp2789) | (tmp2776 & tmp2789);
  wire tmp2791;
  assign tmp2791 = (tmp2710 & tmp2750) | (tmp2710 & tmp2790) | (tmp2750 & tmp2790);
  wire tmp2792;
  assign tmp2792 = 1'b0;
  wire tmp2793;
  assign tmp2793 = 1'b0;
  wire tmp2794;
  assign tmp2794 = 1'b0;
  wire tmp2795;
  assign tmp2795 = (tmp2792 & tmp2793) | (tmp2792 & tmp2794) | (tmp2793 & tmp2794);
  wire tmp2796;
  assign tmp2796 = 1'b0;
  wire tmp2797;
  assign tmp2797 = 1'b0;
  wire tmp2798;
  assign tmp2798 = 1'b0;
  wire tmp2799;
  assign tmp2799 = (tmp2796 & tmp2797) | (tmp2796 & tmp2798) | (tmp2797 & tmp2798);
  wire tmp2800;
  assign tmp2800 = 1'b0;
  wire tmp2801;
  assign tmp2801 = 1'b0;
  wire tmp2802;
  assign tmp2802 = 1'b0;
  wire tmp2803;
  assign tmp2803 = (tmp2800 & tmp2801) | (tmp2800 & tmp2802) | (tmp2801 & tmp2802);
  wire tmp2804;
  assign tmp2804 = (tmp2795 & tmp2799) | (tmp2795 & tmp2803) | (tmp2799 & tmp2803);
  wire tmp2805;
  assign tmp2805 = 1'b0;
  wire tmp2806;
  assign tmp2806 = 1'b0;
  wire tmp2807;
  assign tmp2807 = 1'b0;
  wire tmp2808;
  assign tmp2808 = (tmp2805 & tmp2806) | (tmp2805 & tmp2807) | (tmp2806 & tmp2807);
  wire tmp2809;
  assign tmp2809 = 1'b0;
  wire tmp2810;
  assign tmp2810 = 1'b1;
  wire tmp2811;
  assign tmp2811 = 1'b0;
  wire tmp2812;
  assign tmp2812 = (tmp2809 & tmp2810) | (tmp2809 & tmp2811) | (tmp2810 & tmp2811);
  wire tmp2813;
  assign tmp2813 = 1'b0;
  wire tmp2814;
  assign tmp2814 = 1'b0;
  wire tmp2815;
  assign tmp2815 = 1'b0;
  wire tmp2816;
  assign tmp2816 = (tmp2813 & tmp2814) | (tmp2813 & tmp2815) | (tmp2814 & tmp2815);
  wire tmp2817;
  assign tmp2817 = (tmp2808 & tmp2812) | (tmp2808 & tmp2816) | (tmp2812 & tmp2816);
  wire tmp2818;
  assign tmp2818 = 1'b0;
  wire tmp2819;
  assign tmp2819 = 1'b0;
  wire tmp2820;
  assign tmp2820 = 1'b0;
  wire tmp2821;
  assign tmp2821 = (tmp2818 & tmp2819) | (tmp2818 & tmp2820) | (tmp2819 & tmp2820);
  wire tmp2822;
  assign tmp2822 = 1'b0;
  wire tmp2823;
  assign tmp2823 = 1'b0;
  wire tmp2824;
  assign tmp2824 = 1'b0;
  wire tmp2825;
  assign tmp2825 = (tmp2822 & tmp2823) | (tmp2822 & tmp2824) | (tmp2823 & tmp2824);
  wire tmp2826;
  assign tmp2826 = 1'b0;
  wire tmp2827;
  assign tmp2827 = 1'b0;
  wire tmp2828;
  assign tmp2828 = 1'b0;
  wire tmp2829;
  assign tmp2829 = (tmp2826 & tmp2827) | (tmp2826 & tmp2828) | (tmp2827 & tmp2828);
  wire tmp2830;
  assign tmp2830 = (tmp2821 & tmp2825) | (tmp2821 & tmp2829) | (tmp2825 & tmp2829);
  wire tmp2831;
  assign tmp2831 = (tmp2804 & tmp2817) | (tmp2804 & tmp2830) | (tmp2817 & tmp2830);
  wire tmp2832;
  assign tmp2832 = 1'b0;
  wire tmp2833;
  assign tmp2833 = 1'b0;
  wire tmp2834;
  assign tmp2834 = 1'b0;
  wire tmp2835;
  assign tmp2835 = (tmp2832 & tmp2833) | (tmp2832 & tmp2834) | (tmp2833 & tmp2834);
  wire tmp2836;
  assign tmp2836 = 1'b0;
  wire tmp2837;
  assign tmp2837 = 1'b1;
  wire tmp2838;
  assign tmp2838 = 1'b0;
  wire tmp2839;
  assign tmp2839 = (tmp2836 & tmp2837) | (tmp2836 & tmp2838) | (tmp2837 & tmp2838);
  wire tmp2840;
  assign tmp2840 = 1'b0;
  wire tmp2841;
  assign tmp2841 = 1'b0;
  wire tmp2842;
  assign tmp2842 = 1'b0;
  wire tmp2843;
  assign tmp2843 = (tmp2840 & tmp2841) | (tmp2840 & tmp2842) | (tmp2841 & tmp2842);
  wire tmp2844;
  assign tmp2844 = (tmp2835 & tmp2839) | (tmp2835 & tmp2843) | (tmp2839 & tmp2843);
  wire tmp2845;
  assign tmp2845 = 1'b0;
  wire tmp2846;
  assign tmp2846 = 1'b1;
  wire tmp2847;
  assign tmp2847 = 1'b0;
  wire tmp2848;
  assign tmp2848 = (tmp2845 & tmp2846) | (tmp2845 & tmp2847) | (tmp2846 & tmp2847);
  wire tmp2849;
  assign tmp2849 = 1'b1;
  wire tmp2850;
  assign tmp2850 = ~pi6;
  wire tmp2851;
  assign tmp2851 = ~pi7;
  wire tmp2852;
  assign tmp2852 = (tmp2849 & tmp2850) | (tmp2849 & tmp2851) | (tmp2850 & tmp2851);
  wire tmp2853;
  assign tmp2853 = 1'b0;
  wire tmp2854;
  assign tmp2854 = ~pi7;
  wire tmp2855;
  assign tmp2855 = 1'b0;
  wire tmp2856;
  assign tmp2856 = (tmp2853 & tmp2854) | (tmp2853 & tmp2855) | (tmp2854 & tmp2855);
  wire tmp2857;
  assign tmp2857 = (tmp2848 & tmp2852) | (tmp2848 & tmp2856) | (tmp2852 & tmp2856);
  wire tmp2858;
  assign tmp2858 = 1'b0;
  wire tmp2859;
  assign tmp2859 = 1'b0;
  wire tmp2860;
  assign tmp2860 = 1'b0;
  wire tmp2861;
  assign tmp2861 = (tmp2858 & tmp2859) | (tmp2858 & tmp2860) | (tmp2859 & tmp2860);
  wire tmp2862;
  assign tmp2862 = 1'b0;
  wire tmp2863;
  assign tmp2863 = ~pi7;
  wire tmp2864;
  assign tmp2864 = 1'b0;
  wire tmp2865;
  assign tmp2865 = (tmp2862 & tmp2863) | (tmp2862 & tmp2864) | (tmp2863 & tmp2864);
  wire tmp2866;
  assign tmp2866 = 1'b0;
  wire tmp2867;
  assign tmp2867 = 1'b0;
  wire tmp2868;
  assign tmp2868 = 1'b0;
  wire tmp2869;
  assign tmp2869 = (tmp2866 & tmp2867) | (tmp2866 & tmp2868) | (tmp2867 & tmp2868);
  wire tmp2870;
  assign tmp2870 = (tmp2861 & tmp2865) | (tmp2861 & tmp2869) | (tmp2865 & tmp2869);
  wire tmp2871;
  assign tmp2871 = (tmp2844 & tmp2857) | (tmp2844 & tmp2870) | (tmp2857 & tmp2870);
  wire tmp2872;
  assign tmp2872 = 1'b0;
  wire tmp2873;
  assign tmp2873 = 1'b0;
  wire tmp2874;
  assign tmp2874 = 1'b0;
  wire tmp2875;
  assign tmp2875 = (tmp2872 & tmp2873) | (tmp2872 & tmp2874) | (tmp2873 & tmp2874);
  wire tmp2876;
  assign tmp2876 = 1'b0;
  wire tmp2877;
  assign tmp2877 = 1'b0;
  wire tmp2878;
  assign tmp2878 = 1'b0;
  wire tmp2879;
  assign tmp2879 = (tmp2876 & tmp2877) | (tmp2876 & tmp2878) | (tmp2877 & tmp2878);
  wire tmp2880;
  assign tmp2880 = 1'b0;
  wire tmp2881;
  assign tmp2881 = 1'b0;
  wire tmp2882;
  assign tmp2882 = 1'b0;
  wire tmp2883;
  assign tmp2883 = (tmp2880 & tmp2881) | (tmp2880 & tmp2882) | (tmp2881 & tmp2882);
  wire tmp2884;
  assign tmp2884 = (tmp2875 & tmp2879) | (tmp2875 & tmp2883) | (tmp2879 & tmp2883);
  wire tmp2885;
  assign tmp2885 = 1'b0;
  wire tmp2886;
  assign tmp2886 = 1'b0;
  wire tmp2887;
  assign tmp2887 = 1'b0;
  wire tmp2888;
  assign tmp2888 = (tmp2885 & tmp2886) | (tmp2885 & tmp2887) | (tmp2886 & tmp2887);
  wire tmp2889;
  assign tmp2889 = 1'b0;
  wire tmp2890;
  assign tmp2890 = ~pi7;
  wire tmp2891;
  assign tmp2891 = 1'b0;
  wire tmp2892;
  assign tmp2892 = (tmp2889 & tmp2890) | (tmp2889 & tmp2891) | (tmp2890 & tmp2891);
  wire tmp2893;
  assign tmp2893 = 1'b0;
  wire tmp2894;
  assign tmp2894 = 1'b0;
  wire tmp2895;
  assign tmp2895 = 1'b0;
  wire tmp2896;
  assign tmp2896 = (tmp2893 & tmp2894) | (tmp2893 & tmp2895) | (tmp2894 & tmp2895);
  wire tmp2897;
  assign tmp2897 = (tmp2888 & tmp2892) | (tmp2888 & tmp2896) | (tmp2892 & tmp2896);
  wire tmp2898;
  assign tmp2898 = 1'b0;
  wire tmp2899;
  assign tmp2899 = 1'b0;
  wire tmp2900;
  assign tmp2900 = 1'b0;
  wire tmp2901;
  assign tmp2901 = (tmp2898 & tmp2899) | (tmp2898 & tmp2900) | (tmp2899 & tmp2900);
  wire tmp2902;
  assign tmp2902 = 1'b0;
  wire tmp2903;
  assign tmp2903 = 1'b0;
  wire tmp2904;
  assign tmp2904 = 1'b0;
  wire tmp2905;
  assign tmp2905 = (tmp2902 & tmp2903) | (tmp2902 & tmp2904) | (tmp2903 & tmp2904);
  wire tmp2906;
  assign tmp2906 = 1'b0;
  wire tmp2907;
  assign tmp2907 = 1'b0;
  wire tmp2908;
  assign tmp2908 = 1'b0;
  wire tmp2909;
  assign tmp2909 = (tmp2906 & tmp2907) | (tmp2906 & tmp2908) | (tmp2907 & tmp2908);
  wire tmp2910;
  assign tmp2910 = (tmp2901 & tmp2905) | (tmp2901 & tmp2909) | (tmp2905 & tmp2909);
  wire tmp2911;
  assign tmp2911 = (tmp2884 & tmp2897) | (tmp2884 & tmp2910) | (tmp2897 & tmp2910);
  wire tmp2912;
  assign tmp2912 = (tmp2831 & tmp2871) | (tmp2831 & tmp2911) | (tmp2871 & tmp2911);
  wire tmp2913;
  assign tmp2913 = (tmp2670 & tmp2791) | (tmp2670 & tmp2912) | (tmp2791 & tmp2912);
  wire tmp2914;
  assign tmp2914 = 1'b0;
  wire tmp2915;
  assign tmp2915 = 1'b0;
  wire tmp2916;
  assign tmp2916 = 1'b0;
  wire tmp2917;
  assign tmp2917 = (tmp2914 & tmp2915) | (tmp2914 & tmp2916) | (tmp2915 & tmp2916);
  wire tmp2918;
  assign tmp2918 = 1'b0;
  wire tmp2919;
  assign tmp2919 = 1'b0;
  wire tmp2920;
  assign tmp2920 = 1'b0;
  wire tmp2921;
  assign tmp2921 = (tmp2918 & tmp2919) | (tmp2918 & tmp2920) | (tmp2919 & tmp2920);
  wire tmp2922;
  assign tmp2922 = 1'b0;
  wire tmp2923;
  assign tmp2923 = 1'b0;
  wire tmp2924;
  assign tmp2924 = 1'b0;
  wire tmp2925;
  assign tmp2925 = (tmp2922 & tmp2923) | (tmp2922 & tmp2924) | (tmp2923 & tmp2924);
  wire tmp2926;
  assign tmp2926 = (tmp2917 & tmp2921) | (tmp2917 & tmp2925) | (tmp2921 & tmp2925);
  wire tmp2927;
  assign tmp2927 = 1'b0;
  wire tmp2928;
  assign tmp2928 = 1'b0;
  wire tmp2929;
  assign tmp2929 = 1'b0;
  wire tmp2930;
  assign tmp2930 = (tmp2927 & tmp2928) | (tmp2927 & tmp2929) | (tmp2928 & tmp2929);
  wire tmp2931;
  assign tmp2931 = 1'b0;
  wire tmp2932;
  assign tmp2932 = 1'b0;
  wire tmp2933;
  assign tmp2933 = 1'b0;
  wire tmp2934;
  assign tmp2934 = (tmp2931 & tmp2932) | (tmp2931 & tmp2933) | (tmp2932 & tmp2933);
  wire tmp2935;
  assign tmp2935 = 1'b0;
  wire tmp2936;
  assign tmp2936 = 1'b0;
  wire tmp2937;
  assign tmp2937 = 1'b0;
  wire tmp2938;
  assign tmp2938 = (tmp2935 & tmp2936) | (tmp2935 & tmp2937) | (tmp2936 & tmp2937);
  wire tmp2939;
  assign tmp2939 = (tmp2930 & tmp2934) | (tmp2930 & tmp2938) | (tmp2934 & tmp2938);
  wire tmp2940;
  assign tmp2940 = 1'b0;
  wire tmp2941;
  assign tmp2941 = 1'b0;
  wire tmp2942;
  assign tmp2942 = 1'b0;
  wire tmp2943;
  assign tmp2943 = (tmp2940 & tmp2941) | (tmp2940 & tmp2942) | (tmp2941 & tmp2942);
  wire tmp2944;
  assign tmp2944 = 1'b0;
  wire tmp2945;
  assign tmp2945 = 1'b0;
  wire tmp2946;
  assign tmp2946 = 1'b0;
  wire tmp2947;
  assign tmp2947 = (tmp2944 & tmp2945) | (tmp2944 & tmp2946) | (tmp2945 & tmp2946);
  wire tmp2948;
  assign tmp2948 = 1'b0;
  wire tmp2949;
  assign tmp2949 = 1'b0;
  wire tmp2950;
  assign tmp2950 = 1'b0;
  wire tmp2951;
  assign tmp2951 = (tmp2948 & tmp2949) | (tmp2948 & tmp2950) | (tmp2949 & tmp2950);
  wire tmp2952;
  assign tmp2952 = (tmp2943 & tmp2947) | (tmp2943 & tmp2951) | (tmp2947 & tmp2951);
  wire tmp2953;
  assign tmp2953 = (tmp2926 & tmp2939) | (tmp2926 & tmp2952) | (tmp2939 & tmp2952);
  wire tmp2954;
  assign tmp2954 = 1'b0;
  wire tmp2955;
  assign tmp2955 = 1'b0;
  wire tmp2956;
  assign tmp2956 = 1'b0;
  wire tmp2957;
  assign tmp2957 = (tmp2954 & tmp2955) | (tmp2954 & tmp2956) | (tmp2955 & tmp2956);
  wire tmp2958;
  assign tmp2958 = 1'b0;
  wire tmp2959;
  assign tmp2959 = 1'b0;
  wire tmp2960;
  assign tmp2960 = 1'b0;
  wire tmp2961;
  assign tmp2961 = (tmp2958 & tmp2959) | (tmp2958 & tmp2960) | (tmp2959 & tmp2960);
  wire tmp2962;
  assign tmp2962 = 1'b0;
  wire tmp2963;
  assign tmp2963 = 1'b0;
  wire tmp2964;
  assign tmp2964 = 1'b0;
  wire tmp2965;
  assign tmp2965 = (tmp2962 & tmp2963) | (tmp2962 & tmp2964) | (tmp2963 & tmp2964);
  wire tmp2966;
  assign tmp2966 = (tmp2957 & tmp2961) | (tmp2957 & tmp2965) | (tmp2961 & tmp2965);
  wire tmp2967;
  assign tmp2967 = 1'b0;
  wire tmp2968;
  assign tmp2968 = 1'b0;
  wire tmp2969;
  assign tmp2969 = 1'b0;
  wire tmp2970;
  assign tmp2970 = (tmp2967 & tmp2968) | (tmp2967 & tmp2969) | (tmp2968 & tmp2969);
  wire tmp2971;
  assign tmp2971 = 1'b0;
  wire tmp2972;
  assign tmp2972 = 1'b1;
  wire tmp2973;
  assign tmp2973 = 1'b0;
  wire tmp2974;
  assign tmp2974 = (tmp2971 & tmp2972) | (tmp2971 & tmp2973) | (tmp2972 & tmp2973);
  wire tmp2975;
  assign tmp2975 = 1'b0;
  wire tmp2976;
  assign tmp2976 = 1'b0;
  wire tmp2977;
  assign tmp2977 = 1'b0;
  wire tmp2978;
  assign tmp2978 = (tmp2975 & tmp2976) | (tmp2975 & tmp2977) | (tmp2976 & tmp2977);
  wire tmp2979;
  assign tmp2979 = (tmp2970 & tmp2974) | (tmp2970 & tmp2978) | (tmp2974 & tmp2978);
  wire tmp2980;
  assign tmp2980 = 1'b0;
  wire tmp2981;
  assign tmp2981 = 1'b0;
  wire tmp2982;
  assign tmp2982 = 1'b0;
  wire tmp2983;
  assign tmp2983 = (tmp2980 & tmp2981) | (tmp2980 & tmp2982) | (tmp2981 & tmp2982);
  wire tmp2984;
  assign tmp2984 = 1'b0;
  wire tmp2985;
  assign tmp2985 = 1'b0;
  wire tmp2986;
  assign tmp2986 = 1'b0;
  wire tmp2987;
  assign tmp2987 = (tmp2984 & tmp2985) | (tmp2984 & tmp2986) | (tmp2985 & tmp2986);
  wire tmp2988;
  assign tmp2988 = 1'b0;
  wire tmp2989;
  assign tmp2989 = 1'b0;
  wire tmp2990;
  assign tmp2990 = 1'b0;
  wire tmp2991;
  assign tmp2991 = (tmp2988 & tmp2989) | (tmp2988 & tmp2990) | (tmp2989 & tmp2990);
  wire tmp2992;
  assign tmp2992 = (tmp2983 & tmp2987) | (tmp2983 & tmp2991) | (tmp2987 & tmp2991);
  wire tmp2993;
  assign tmp2993 = (tmp2966 & tmp2979) | (tmp2966 & tmp2992) | (tmp2979 & tmp2992);
  wire tmp2994;
  assign tmp2994 = 1'b0;
  wire tmp2995;
  assign tmp2995 = 1'b0;
  wire tmp2996;
  assign tmp2996 = 1'b0;
  wire tmp2997;
  assign tmp2997 = (tmp2994 & tmp2995) | (tmp2994 & tmp2996) | (tmp2995 & tmp2996);
  wire tmp2998;
  assign tmp2998 = 1'b0;
  wire tmp2999;
  assign tmp2999 = 1'b0;
  wire tmp3000;
  assign tmp3000 = 1'b0;
  wire tmp3001;
  assign tmp3001 = (tmp2998 & tmp2999) | (tmp2998 & tmp3000) | (tmp2999 & tmp3000);
  wire tmp3002;
  assign tmp3002 = 1'b0;
  wire tmp3003;
  assign tmp3003 = 1'b0;
  wire tmp3004;
  assign tmp3004 = 1'b0;
  wire tmp3005;
  assign tmp3005 = (tmp3002 & tmp3003) | (tmp3002 & tmp3004) | (tmp3003 & tmp3004);
  wire tmp3006;
  assign tmp3006 = (tmp2997 & tmp3001) | (tmp2997 & tmp3005) | (tmp3001 & tmp3005);
  wire tmp3007;
  assign tmp3007 = 1'b0;
  wire tmp3008;
  assign tmp3008 = 1'b0;
  wire tmp3009;
  assign tmp3009 = 1'b0;
  wire tmp3010;
  assign tmp3010 = (tmp3007 & tmp3008) | (tmp3007 & tmp3009) | (tmp3008 & tmp3009);
  wire tmp3011;
  assign tmp3011 = 1'b0;
  wire tmp3012;
  assign tmp3012 = 1'b0;
  wire tmp3013;
  assign tmp3013 = 1'b0;
  wire tmp3014;
  assign tmp3014 = (tmp3011 & tmp3012) | (tmp3011 & tmp3013) | (tmp3012 & tmp3013);
  wire tmp3015;
  assign tmp3015 = 1'b0;
  wire tmp3016;
  assign tmp3016 = 1'b0;
  wire tmp3017;
  assign tmp3017 = 1'b0;
  wire tmp3018;
  assign tmp3018 = (tmp3015 & tmp3016) | (tmp3015 & tmp3017) | (tmp3016 & tmp3017);
  wire tmp3019;
  assign tmp3019 = (tmp3010 & tmp3014) | (tmp3010 & tmp3018) | (tmp3014 & tmp3018);
  wire tmp3020;
  assign tmp3020 = 1'b0;
  wire tmp3021;
  assign tmp3021 = 1'b0;
  wire tmp3022;
  assign tmp3022 = 1'b0;
  wire tmp3023;
  assign tmp3023 = (tmp3020 & tmp3021) | (tmp3020 & tmp3022) | (tmp3021 & tmp3022);
  wire tmp3024;
  assign tmp3024 = 1'b0;
  wire tmp3025;
  assign tmp3025 = 1'b0;
  wire tmp3026;
  assign tmp3026 = 1'b0;
  wire tmp3027;
  assign tmp3027 = (tmp3024 & tmp3025) | (tmp3024 & tmp3026) | (tmp3025 & tmp3026);
  wire tmp3028;
  assign tmp3028 = 1'b0;
  wire tmp3029;
  assign tmp3029 = 1'b0;
  wire tmp3030;
  assign tmp3030 = 1'b0;
  wire tmp3031;
  assign tmp3031 = (tmp3028 & tmp3029) | (tmp3028 & tmp3030) | (tmp3029 & tmp3030);
  wire tmp3032;
  assign tmp3032 = (tmp3023 & tmp3027) | (tmp3023 & tmp3031) | (tmp3027 & tmp3031);
  wire tmp3033;
  assign tmp3033 = (tmp3006 & tmp3019) | (tmp3006 & tmp3032) | (tmp3019 & tmp3032);
  wire tmp3034;
  assign tmp3034 = (tmp2953 & tmp2993) | (tmp2953 & tmp3033) | (tmp2993 & tmp3033);
  wire tmp3035;
  assign tmp3035 = 1'b0;
  wire tmp3036;
  assign tmp3036 = 1'b0;
  wire tmp3037;
  assign tmp3037 = 1'b0;
  wire tmp3038;
  assign tmp3038 = (tmp3035 & tmp3036) | (tmp3035 & tmp3037) | (tmp3036 & tmp3037);
  wire tmp3039;
  assign tmp3039 = 1'b0;
  wire tmp3040;
  assign tmp3040 = 1'b0;
  wire tmp3041;
  assign tmp3041 = 1'b0;
  wire tmp3042;
  assign tmp3042 = (tmp3039 & tmp3040) | (tmp3039 & tmp3041) | (tmp3040 & tmp3041);
  wire tmp3043;
  assign tmp3043 = 1'b0;
  wire tmp3044;
  assign tmp3044 = 1'b0;
  wire tmp3045;
  assign tmp3045 = 1'b0;
  wire tmp3046;
  assign tmp3046 = (tmp3043 & tmp3044) | (tmp3043 & tmp3045) | (tmp3044 & tmp3045);
  wire tmp3047;
  assign tmp3047 = (tmp3038 & tmp3042) | (tmp3038 & tmp3046) | (tmp3042 & tmp3046);
  wire tmp3048;
  assign tmp3048 = 1'b0;
  wire tmp3049;
  assign tmp3049 = 1'b0;
  wire tmp3050;
  assign tmp3050 = 1'b0;
  wire tmp3051;
  assign tmp3051 = (tmp3048 & tmp3049) | (tmp3048 & tmp3050) | (tmp3049 & tmp3050);
  wire tmp3052;
  assign tmp3052 = 1'b0;
  wire tmp3053;
  assign tmp3053 = 1'b1;
  wire tmp3054;
  assign tmp3054 = 1'b0;
  wire tmp3055;
  assign tmp3055 = (tmp3052 & tmp3053) | (tmp3052 & tmp3054) | (tmp3053 & tmp3054);
  wire tmp3056;
  assign tmp3056 = 1'b0;
  wire tmp3057;
  assign tmp3057 = 1'b0;
  wire tmp3058;
  assign tmp3058 = 1'b0;
  wire tmp3059;
  assign tmp3059 = (tmp3056 & tmp3057) | (tmp3056 & tmp3058) | (tmp3057 & tmp3058);
  wire tmp3060;
  assign tmp3060 = (tmp3051 & tmp3055) | (tmp3051 & tmp3059) | (tmp3055 & tmp3059);
  wire tmp3061;
  assign tmp3061 = 1'b0;
  wire tmp3062;
  assign tmp3062 = 1'b0;
  wire tmp3063;
  assign tmp3063 = 1'b0;
  wire tmp3064;
  assign tmp3064 = (tmp3061 & tmp3062) | (tmp3061 & tmp3063) | (tmp3062 & tmp3063);
  wire tmp3065;
  assign tmp3065 = 1'b0;
  wire tmp3066;
  assign tmp3066 = 1'b0;
  wire tmp3067;
  assign tmp3067 = 1'b0;
  wire tmp3068;
  assign tmp3068 = (tmp3065 & tmp3066) | (tmp3065 & tmp3067) | (tmp3066 & tmp3067);
  wire tmp3069;
  assign tmp3069 = 1'b0;
  wire tmp3070;
  assign tmp3070 = 1'b0;
  wire tmp3071;
  assign tmp3071 = 1'b0;
  wire tmp3072;
  assign tmp3072 = (tmp3069 & tmp3070) | (tmp3069 & tmp3071) | (tmp3070 & tmp3071);
  wire tmp3073;
  assign tmp3073 = (tmp3064 & tmp3068) | (tmp3064 & tmp3072) | (tmp3068 & tmp3072);
  wire tmp3074;
  assign tmp3074 = (tmp3047 & tmp3060) | (tmp3047 & tmp3073) | (tmp3060 & tmp3073);
  wire tmp3075;
  assign tmp3075 = 1'b0;
  wire tmp3076;
  assign tmp3076 = 1'b0;
  wire tmp3077;
  assign tmp3077 = 1'b0;
  wire tmp3078;
  assign tmp3078 = (tmp3075 & tmp3076) | (tmp3075 & tmp3077) | (tmp3076 & tmp3077);
  wire tmp3079;
  assign tmp3079 = 1'b0;
  wire tmp3080;
  assign tmp3080 = 1'b1;
  wire tmp3081;
  assign tmp3081 = 1'b0;
  wire tmp3082;
  assign tmp3082 = (tmp3079 & tmp3080) | (tmp3079 & tmp3081) | (tmp3080 & tmp3081);
  wire tmp3083;
  assign tmp3083 = 1'b0;
  wire tmp3084;
  assign tmp3084 = 1'b0;
  wire tmp3085;
  assign tmp3085 = 1'b0;
  wire tmp3086;
  assign tmp3086 = (tmp3083 & tmp3084) | (tmp3083 & tmp3085) | (tmp3084 & tmp3085);
  wire tmp3087;
  assign tmp3087 = (tmp3078 & tmp3082) | (tmp3078 & tmp3086) | (tmp3082 & tmp3086);
  wire tmp3088;
  assign tmp3088 = 1'b0;
  wire tmp3089;
  assign tmp3089 = 1'b1;
  wire tmp3090;
  assign tmp3090 = 1'b0;
  wire tmp3091;
  assign tmp3091 = (tmp3088 & tmp3089) | (tmp3088 & tmp3090) | (tmp3089 & tmp3090);
  wire tmp3092;
  assign tmp3092 = 1'b1;
  wire tmp3093;
  assign tmp3093 = ~pi6;
  wire tmp3094;
  assign tmp3094 = ~pi7;
  wire tmp3095;
  assign tmp3095 = (tmp3092 & tmp3093) | (tmp3092 & tmp3094) | (tmp3093 & tmp3094);
  wire tmp3096;
  assign tmp3096 = 1'b0;
  wire tmp3097;
  assign tmp3097 = ~pi7;
  wire tmp3098;
  assign tmp3098 = 1'b0;
  wire tmp3099;
  assign tmp3099 = (tmp3096 & tmp3097) | (tmp3096 & tmp3098) | (tmp3097 & tmp3098);
  wire tmp3100;
  assign tmp3100 = (tmp3091 & tmp3095) | (tmp3091 & tmp3099) | (tmp3095 & tmp3099);
  wire tmp3101;
  assign tmp3101 = 1'b0;
  wire tmp3102;
  assign tmp3102 = 1'b0;
  wire tmp3103;
  assign tmp3103 = 1'b0;
  wire tmp3104;
  assign tmp3104 = (tmp3101 & tmp3102) | (tmp3101 & tmp3103) | (tmp3102 & tmp3103);
  wire tmp3105;
  assign tmp3105 = 1'b0;
  wire tmp3106;
  assign tmp3106 = ~pi7;
  wire tmp3107;
  assign tmp3107 = 1'b0;
  wire tmp3108;
  assign tmp3108 = (tmp3105 & tmp3106) | (tmp3105 & tmp3107) | (tmp3106 & tmp3107);
  wire tmp3109;
  assign tmp3109 = 1'b0;
  wire tmp3110;
  assign tmp3110 = 1'b0;
  wire tmp3111;
  assign tmp3111 = 1'b0;
  wire tmp3112;
  assign tmp3112 = (tmp3109 & tmp3110) | (tmp3109 & tmp3111) | (tmp3110 & tmp3111);
  wire tmp3113;
  assign tmp3113 = (tmp3104 & tmp3108) | (tmp3104 & tmp3112) | (tmp3108 & tmp3112);
  wire tmp3114;
  assign tmp3114 = (tmp3087 & tmp3100) | (tmp3087 & tmp3113) | (tmp3100 & tmp3113);
  wire tmp3115;
  assign tmp3115 = 1'b0;
  wire tmp3116;
  assign tmp3116 = 1'b0;
  wire tmp3117;
  assign tmp3117 = 1'b0;
  wire tmp3118;
  assign tmp3118 = (tmp3115 & tmp3116) | (tmp3115 & tmp3117) | (tmp3116 & tmp3117);
  wire tmp3119;
  assign tmp3119 = 1'b0;
  wire tmp3120;
  assign tmp3120 = 1'b0;
  wire tmp3121;
  assign tmp3121 = 1'b0;
  wire tmp3122;
  assign tmp3122 = (tmp3119 & tmp3120) | (tmp3119 & tmp3121) | (tmp3120 & tmp3121);
  wire tmp3123;
  assign tmp3123 = 1'b0;
  wire tmp3124;
  assign tmp3124 = 1'b0;
  wire tmp3125;
  assign tmp3125 = 1'b0;
  wire tmp3126;
  assign tmp3126 = (tmp3123 & tmp3124) | (tmp3123 & tmp3125) | (tmp3124 & tmp3125);
  wire tmp3127;
  assign tmp3127 = (tmp3118 & tmp3122) | (tmp3118 & tmp3126) | (tmp3122 & tmp3126);
  wire tmp3128;
  assign tmp3128 = 1'b0;
  wire tmp3129;
  assign tmp3129 = 1'b0;
  wire tmp3130;
  assign tmp3130 = 1'b0;
  wire tmp3131;
  assign tmp3131 = (tmp3128 & tmp3129) | (tmp3128 & tmp3130) | (tmp3129 & tmp3130);
  wire tmp3132;
  assign tmp3132 = 1'b0;
  wire tmp3133;
  assign tmp3133 = ~pi7;
  wire tmp3134;
  assign tmp3134 = 1'b0;
  wire tmp3135;
  assign tmp3135 = (tmp3132 & tmp3133) | (tmp3132 & tmp3134) | (tmp3133 & tmp3134);
  wire tmp3136;
  assign tmp3136 = 1'b0;
  wire tmp3137;
  assign tmp3137 = 1'b0;
  wire tmp3138;
  assign tmp3138 = 1'b0;
  wire tmp3139;
  assign tmp3139 = (tmp3136 & tmp3137) | (tmp3136 & tmp3138) | (tmp3137 & tmp3138);
  wire tmp3140;
  assign tmp3140 = (tmp3131 & tmp3135) | (tmp3131 & tmp3139) | (tmp3135 & tmp3139);
  wire tmp3141;
  assign tmp3141 = 1'b0;
  wire tmp3142;
  assign tmp3142 = 1'b0;
  wire tmp3143;
  assign tmp3143 = 1'b0;
  wire tmp3144;
  assign tmp3144 = (tmp3141 & tmp3142) | (tmp3141 & tmp3143) | (tmp3142 & tmp3143);
  wire tmp3145;
  assign tmp3145 = 1'b0;
  wire tmp3146;
  assign tmp3146 = 1'b0;
  wire tmp3147;
  assign tmp3147 = 1'b0;
  wire tmp3148;
  assign tmp3148 = (tmp3145 & tmp3146) | (tmp3145 & tmp3147) | (tmp3146 & tmp3147);
  wire tmp3149;
  assign tmp3149 = 1'b0;
  wire tmp3150;
  assign tmp3150 = 1'b0;
  wire tmp3151;
  assign tmp3151 = 1'b0;
  wire tmp3152;
  assign tmp3152 = (tmp3149 & tmp3150) | (tmp3149 & tmp3151) | (tmp3150 & tmp3151);
  wire tmp3153;
  assign tmp3153 = (tmp3144 & tmp3148) | (tmp3144 & tmp3152) | (tmp3148 & tmp3152);
  wire tmp3154;
  assign tmp3154 = (tmp3127 & tmp3140) | (tmp3127 & tmp3153) | (tmp3140 & tmp3153);
  wire tmp3155;
  assign tmp3155 = (tmp3074 & tmp3114) | (tmp3074 & tmp3154) | (tmp3114 & tmp3154);
  wire tmp3156;
  assign tmp3156 = 1'b0;
  wire tmp3157;
  assign tmp3157 = 1'b0;
  wire tmp3158;
  assign tmp3158 = 1'b0;
  wire tmp3159;
  assign tmp3159 = (tmp3156 & tmp3157) | (tmp3156 & tmp3158) | (tmp3157 & tmp3158);
  wire tmp3160;
  assign tmp3160 = 1'b0;
  wire tmp3161;
  assign tmp3161 = 1'b0;
  wire tmp3162;
  assign tmp3162 = 1'b0;
  wire tmp3163;
  assign tmp3163 = (tmp3160 & tmp3161) | (tmp3160 & tmp3162) | (tmp3161 & tmp3162);
  wire tmp3164;
  assign tmp3164 = 1'b0;
  wire tmp3165;
  assign tmp3165 = 1'b0;
  wire tmp3166;
  assign tmp3166 = 1'b0;
  wire tmp3167;
  assign tmp3167 = (tmp3164 & tmp3165) | (tmp3164 & tmp3166) | (tmp3165 & tmp3166);
  wire tmp3168;
  assign tmp3168 = (tmp3159 & tmp3163) | (tmp3159 & tmp3167) | (tmp3163 & tmp3167);
  wire tmp3169;
  assign tmp3169 = 1'b0;
  wire tmp3170;
  assign tmp3170 = 1'b0;
  wire tmp3171;
  assign tmp3171 = 1'b0;
  wire tmp3172;
  assign tmp3172 = (tmp3169 & tmp3170) | (tmp3169 & tmp3171) | (tmp3170 & tmp3171);
  wire tmp3173;
  assign tmp3173 = 1'b0;
  wire tmp3174;
  assign tmp3174 = 1'b0;
  wire tmp3175;
  assign tmp3175 = 1'b0;
  wire tmp3176;
  assign tmp3176 = (tmp3173 & tmp3174) | (tmp3173 & tmp3175) | (tmp3174 & tmp3175);
  wire tmp3177;
  assign tmp3177 = 1'b0;
  wire tmp3178;
  assign tmp3178 = 1'b0;
  wire tmp3179;
  assign tmp3179 = 1'b0;
  wire tmp3180;
  assign tmp3180 = (tmp3177 & tmp3178) | (tmp3177 & tmp3179) | (tmp3178 & tmp3179);
  wire tmp3181;
  assign tmp3181 = (tmp3172 & tmp3176) | (tmp3172 & tmp3180) | (tmp3176 & tmp3180);
  wire tmp3182;
  assign tmp3182 = 1'b0;
  wire tmp3183;
  assign tmp3183 = 1'b0;
  wire tmp3184;
  assign tmp3184 = 1'b0;
  wire tmp3185;
  assign tmp3185 = (tmp3182 & tmp3183) | (tmp3182 & tmp3184) | (tmp3183 & tmp3184);
  wire tmp3186;
  assign tmp3186 = 1'b0;
  wire tmp3187;
  assign tmp3187 = 1'b0;
  wire tmp3188;
  assign tmp3188 = 1'b0;
  wire tmp3189;
  assign tmp3189 = (tmp3186 & tmp3187) | (tmp3186 & tmp3188) | (tmp3187 & tmp3188);
  wire tmp3190;
  assign tmp3190 = 1'b0;
  wire tmp3191;
  assign tmp3191 = 1'b0;
  wire tmp3192;
  assign tmp3192 = 1'b0;
  wire tmp3193;
  assign tmp3193 = (tmp3190 & tmp3191) | (tmp3190 & tmp3192) | (tmp3191 & tmp3192);
  wire tmp3194;
  assign tmp3194 = (tmp3185 & tmp3189) | (tmp3185 & tmp3193) | (tmp3189 & tmp3193);
  wire tmp3195;
  assign tmp3195 = (tmp3168 & tmp3181) | (tmp3168 & tmp3194) | (tmp3181 & tmp3194);
  wire tmp3196;
  assign tmp3196 = 1'b0;
  wire tmp3197;
  assign tmp3197 = 1'b0;
  wire tmp3198;
  assign tmp3198 = 1'b0;
  wire tmp3199;
  assign tmp3199 = (tmp3196 & tmp3197) | (tmp3196 & tmp3198) | (tmp3197 & tmp3198);
  wire tmp3200;
  assign tmp3200 = 1'b0;
  wire tmp3201;
  assign tmp3201 = 1'b0;
  wire tmp3202;
  assign tmp3202 = 1'b0;
  wire tmp3203;
  assign tmp3203 = (tmp3200 & tmp3201) | (tmp3200 & tmp3202) | (tmp3201 & tmp3202);
  wire tmp3204;
  assign tmp3204 = 1'b0;
  wire tmp3205;
  assign tmp3205 = 1'b0;
  wire tmp3206;
  assign tmp3206 = 1'b0;
  wire tmp3207;
  assign tmp3207 = (tmp3204 & tmp3205) | (tmp3204 & tmp3206) | (tmp3205 & tmp3206);
  wire tmp3208;
  assign tmp3208 = (tmp3199 & tmp3203) | (tmp3199 & tmp3207) | (tmp3203 & tmp3207);
  wire tmp3209;
  assign tmp3209 = 1'b0;
  wire tmp3210;
  assign tmp3210 = 1'b0;
  wire tmp3211;
  assign tmp3211 = 1'b0;
  wire tmp3212;
  assign tmp3212 = (tmp3209 & tmp3210) | (tmp3209 & tmp3211) | (tmp3210 & tmp3211);
  wire tmp3213;
  assign tmp3213 = 1'b0;
  wire tmp3214;
  assign tmp3214 = ~pi7;
  wire tmp3215;
  assign tmp3215 = 1'b0;
  wire tmp3216;
  assign tmp3216 = (tmp3213 & tmp3214) | (tmp3213 & tmp3215) | (tmp3214 & tmp3215);
  wire tmp3217;
  assign tmp3217 = 1'b0;
  wire tmp3218;
  assign tmp3218 = 1'b0;
  wire tmp3219;
  assign tmp3219 = 1'b0;
  wire tmp3220;
  assign tmp3220 = (tmp3217 & tmp3218) | (tmp3217 & tmp3219) | (tmp3218 & tmp3219);
  wire tmp3221;
  assign tmp3221 = (tmp3212 & tmp3216) | (tmp3212 & tmp3220) | (tmp3216 & tmp3220);
  wire tmp3222;
  assign tmp3222 = 1'b0;
  wire tmp3223;
  assign tmp3223 = 1'b0;
  wire tmp3224;
  assign tmp3224 = 1'b0;
  wire tmp3225;
  assign tmp3225 = (tmp3222 & tmp3223) | (tmp3222 & tmp3224) | (tmp3223 & tmp3224);
  wire tmp3226;
  assign tmp3226 = 1'b0;
  wire tmp3227;
  assign tmp3227 = 1'b0;
  wire tmp3228;
  assign tmp3228 = 1'b0;
  wire tmp3229;
  assign tmp3229 = (tmp3226 & tmp3227) | (tmp3226 & tmp3228) | (tmp3227 & tmp3228);
  wire tmp3230;
  assign tmp3230 = 1'b0;
  wire tmp3231;
  assign tmp3231 = 1'b0;
  wire tmp3232;
  assign tmp3232 = 1'b0;
  wire tmp3233;
  assign tmp3233 = (tmp3230 & tmp3231) | (tmp3230 & tmp3232) | (tmp3231 & tmp3232);
  wire tmp3234;
  assign tmp3234 = (tmp3225 & tmp3229) | (tmp3225 & tmp3233) | (tmp3229 & tmp3233);
  wire tmp3235;
  assign tmp3235 = (tmp3208 & tmp3221) | (tmp3208 & tmp3234) | (tmp3221 & tmp3234);
  wire tmp3236;
  assign tmp3236 = 1'b0;
  wire tmp3237;
  assign tmp3237 = 1'b0;
  wire tmp3238;
  assign tmp3238 = 1'b0;
  wire tmp3239;
  assign tmp3239 = (tmp3236 & tmp3237) | (tmp3236 & tmp3238) | (tmp3237 & tmp3238);
  wire tmp3240;
  assign tmp3240 = 1'b0;
  wire tmp3241;
  assign tmp3241 = 1'b0;
  wire tmp3242;
  assign tmp3242 = 1'b0;
  wire tmp3243;
  assign tmp3243 = (tmp3240 & tmp3241) | (tmp3240 & tmp3242) | (tmp3241 & tmp3242);
  wire tmp3244;
  assign tmp3244 = 1'b0;
  wire tmp3245;
  assign tmp3245 = 1'b0;
  wire tmp3246;
  assign tmp3246 = 1'b0;
  wire tmp3247;
  assign tmp3247 = (tmp3244 & tmp3245) | (tmp3244 & tmp3246) | (tmp3245 & tmp3246);
  wire tmp3248;
  assign tmp3248 = (tmp3239 & tmp3243) | (tmp3239 & tmp3247) | (tmp3243 & tmp3247);
  wire tmp3249;
  assign tmp3249 = 1'b0;
  wire tmp3250;
  assign tmp3250 = 1'b0;
  wire tmp3251;
  assign tmp3251 = 1'b0;
  wire tmp3252;
  assign tmp3252 = (tmp3249 & tmp3250) | (tmp3249 & tmp3251) | (tmp3250 & tmp3251);
  wire tmp3253;
  assign tmp3253 = 1'b0;
  wire tmp3254;
  assign tmp3254 = 1'b0;
  wire tmp3255;
  assign tmp3255 = 1'b0;
  wire tmp3256;
  assign tmp3256 = (tmp3253 & tmp3254) | (tmp3253 & tmp3255) | (tmp3254 & tmp3255);
  wire tmp3257;
  assign tmp3257 = 1'b0;
  wire tmp3258;
  assign tmp3258 = 1'b0;
  wire tmp3259;
  assign tmp3259 = 1'b0;
  wire tmp3260;
  assign tmp3260 = (tmp3257 & tmp3258) | (tmp3257 & tmp3259) | (tmp3258 & tmp3259);
  wire tmp3261;
  assign tmp3261 = (tmp3252 & tmp3256) | (tmp3252 & tmp3260) | (tmp3256 & tmp3260);
  wire tmp3262;
  assign tmp3262 = 1'b0;
  wire tmp3263;
  assign tmp3263 = 1'b0;
  wire tmp3264;
  assign tmp3264 = 1'b0;
  wire tmp3265;
  assign tmp3265 = (tmp3262 & tmp3263) | (tmp3262 & tmp3264) | (tmp3263 & tmp3264);
  wire tmp3266;
  assign tmp3266 = 1'b0;
  wire tmp3267;
  assign tmp3267 = 1'b0;
  wire tmp3268;
  assign tmp3268 = 1'b0;
  wire tmp3269;
  assign tmp3269 = (tmp3266 & tmp3267) | (tmp3266 & tmp3268) | (tmp3267 & tmp3268);
  wire tmp3270;
  assign tmp3270 = 1'b0;
  wire tmp3271;
  assign tmp3271 = 1'b0;
  wire tmp3272;
  assign tmp3272 = 1'b0;
  wire tmp3273;
  assign tmp3273 = (tmp3270 & tmp3271) | (tmp3270 & tmp3272) | (tmp3271 & tmp3272);
  wire tmp3274;
  assign tmp3274 = (tmp3265 & tmp3269) | (tmp3265 & tmp3273) | (tmp3269 & tmp3273);
  wire tmp3275;
  assign tmp3275 = (tmp3248 & tmp3261) | (tmp3248 & tmp3274) | (tmp3261 & tmp3274);
  wire tmp3276;
  assign tmp3276 = (tmp3195 & tmp3235) | (tmp3195 & tmp3275) | (tmp3235 & tmp3275);
  wire tmp3277;
  assign tmp3277 = (tmp3034 & tmp3155) | (tmp3034 & tmp3276) | (tmp3155 & tmp3276);
  wire tmp3278;
  assign tmp3278 = (tmp2549 & tmp2913) | (tmp2549 & tmp3277) | (tmp2913 & tmp3277);
  wire tmp3279;
  assign tmp3279 = (tmp1092 & tmp2185) | (tmp1092 & tmp3278) | (tmp2185 & tmp3278);
  wire tmp3280;
  assign tmp3280 = pi1;
  wire tmp3281;
  assign tmp3281 = pi2;
  wire tmp3282;
  assign tmp3282 = 1'b0;
  wire tmp3283;
  assign tmp3283 = (tmp3280 & tmp3281) | (tmp3280 & tmp3282) | (tmp3281 & tmp3282);
  wire tmp3284;
  assign tmp3284 = pi2;
  wire tmp3285;
  assign tmp3285 = pi3;
  wire tmp3286;
  assign tmp3286 = 1'b0;
  wire tmp3287;
  assign tmp3287 = (tmp3284 & tmp3285) | (tmp3284 & tmp3286) | (tmp3285 & tmp3286);
  wire tmp3288;
  assign tmp3288 = 1'b0;
  wire tmp3289;
  assign tmp3289 = 1'b0;
  wire tmp3290;
  assign tmp3290 = 1'b0;
  wire tmp3291;
  assign tmp3291 = (tmp3288 & tmp3289) | (tmp3288 & tmp3290) | (tmp3289 & tmp3290);
  wire tmp3292;
  assign tmp3292 = (tmp3283 & tmp3287) | (tmp3283 & tmp3291) | (tmp3287 & tmp3291);
  wire tmp3293;
  assign tmp3293 = pi2;
  wire tmp3294;
  assign tmp3294 = pi3;
  wire tmp3295;
  assign tmp3295 = 1'b0;
  wire tmp3296;
  assign tmp3296 = (tmp3293 & tmp3294) | (tmp3293 & tmp3295) | (tmp3294 & tmp3295);
  wire tmp3297;
  assign tmp3297 = pi3;
  wire tmp3298;
  assign tmp3298 = 1'b1;
  wire tmp3299;
  assign tmp3299 = 1'b0;
  wire tmp3300;
  assign tmp3300 = (tmp3297 & tmp3298) | (tmp3297 & tmp3299) | (tmp3298 & tmp3299);
  wire tmp3301;
  assign tmp3301 = 1'b0;
  wire tmp3302;
  assign tmp3302 = 1'b0;
  wire tmp3303;
  assign tmp3303 = 1'b0;
  wire tmp3304;
  assign tmp3304 = (tmp3301 & tmp3302) | (tmp3301 & tmp3303) | (tmp3302 & tmp3303);
  wire tmp3305;
  assign tmp3305 = (tmp3296 & tmp3300) | (tmp3296 & tmp3304) | (tmp3300 & tmp3304);
  wire tmp3306;
  assign tmp3306 = 1'b0;
  wire tmp3307;
  assign tmp3307 = 1'b0;
  wire tmp3308;
  assign tmp3308 = 1'b0;
  wire tmp3309;
  assign tmp3309 = (tmp3306 & tmp3307) | (tmp3306 & tmp3308) | (tmp3307 & tmp3308);
  wire tmp3310;
  assign tmp3310 = 1'b0;
  wire tmp3311;
  assign tmp3311 = 1'b0;
  wire tmp3312;
  assign tmp3312 = 1'b0;
  wire tmp3313;
  assign tmp3313 = (tmp3310 & tmp3311) | (tmp3310 & tmp3312) | (tmp3311 & tmp3312);
  wire tmp3314;
  assign tmp3314 = 1'b0;
  wire tmp3315;
  assign tmp3315 = 1'b0;
  wire tmp3316;
  assign tmp3316 = 1'b0;
  wire tmp3317;
  assign tmp3317 = (tmp3314 & tmp3315) | (tmp3314 & tmp3316) | (tmp3315 & tmp3316);
  wire tmp3318;
  assign tmp3318 = (tmp3309 & tmp3313) | (tmp3309 & tmp3317) | (tmp3313 & tmp3317);
  wire tmp3319;
  assign tmp3319 = (tmp3292 & tmp3305) | (tmp3292 & tmp3318) | (tmp3305 & tmp3318);
  wire tmp3320;
  assign tmp3320 = pi2;
  wire tmp3321;
  assign tmp3321 = pi3;
  wire tmp3322;
  assign tmp3322 = 1'b0;
  wire tmp3323;
  assign tmp3323 = (tmp3320 & tmp3321) | (tmp3320 & tmp3322) | (tmp3321 & tmp3322);
  wire tmp3324;
  assign tmp3324 = pi3;
  wire tmp3325;
  assign tmp3325 = 1'b1;
  wire tmp3326;
  assign tmp3326 = 1'b0;
  wire tmp3327;
  assign tmp3327 = (tmp3324 & tmp3325) | (tmp3324 & tmp3326) | (tmp3325 & tmp3326);
  wire tmp3328;
  assign tmp3328 = 1'b0;
  wire tmp3329;
  assign tmp3329 = 1'b0;
  wire tmp3330;
  assign tmp3330 = 1'b0;
  wire tmp3331;
  assign tmp3331 = (tmp3328 & tmp3329) | (tmp3328 & tmp3330) | (tmp3329 & tmp3330);
  wire tmp3332;
  assign tmp3332 = (tmp3323 & tmp3327) | (tmp3323 & tmp3331) | (tmp3327 & tmp3331);
  wire tmp3333;
  assign tmp3333 = pi3;
  wire tmp3334;
  assign tmp3334 = 1'b1;
  wire tmp3335;
  assign tmp3335 = 1'b0;
  wire tmp3336;
  assign tmp3336 = (tmp3333 & tmp3334) | (tmp3333 & tmp3335) | (tmp3334 & tmp3335);
  wire tmp3337;
  assign tmp3337 = 1'b1;
  wire tmp3338;
  assign tmp3338 = 1'b1;
  wire tmp3339;
  assign tmp3339 = 1'b1;
  wire tmp3340;
  assign tmp3340 = (tmp3337 & tmp3338) | (tmp3337 & tmp3339) | (tmp3338 & tmp3339);
  wire tmp3341;
  assign tmp3341 = 1'b0;
  wire tmp3342;
  assign tmp3342 = 1'b1;
  wire tmp3343;
  assign tmp3343 = 1'b0;
  wire tmp3344;
  assign tmp3344 = (tmp3341 & tmp3342) | (tmp3341 & tmp3343) | (tmp3342 & tmp3343);
  wire tmp3345;
  assign tmp3345 = (tmp3336 & tmp3340) | (tmp3336 & tmp3344) | (tmp3340 & tmp3344);
  wire tmp3346;
  assign tmp3346 = 1'b0;
  wire tmp3347;
  assign tmp3347 = 1'b0;
  wire tmp3348;
  assign tmp3348 = 1'b0;
  wire tmp3349;
  assign tmp3349 = (tmp3346 & tmp3347) | (tmp3346 & tmp3348) | (tmp3347 & tmp3348);
  wire tmp3350;
  assign tmp3350 = 1'b0;
  wire tmp3351;
  assign tmp3351 = 1'b1;
  wire tmp3352;
  assign tmp3352 = 1'b0;
  wire tmp3353;
  assign tmp3353 = (tmp3350 & tmp3351) | (tmp3350 & tmp3352) | (tmp3351 & tmp3352);
  wire tmp3354;
  assign tmp3354 = 1'b0;
  wire tmp3355;
  assign tmp3355 = 1'b0;
  wire tmp3356;
  assign tmp3356 = 1'b0;
  wire tmp3357;
  assign tmp3357 = (tmp3354 & tmp3355) | (tmp3354 & tmp3356) | (tmp3355 & tmp3356);
  wire tmp3358;
  assign tmp3358 = (tmp3349 & tmp3353) | (tmp3349 & tmp3357) | (tmp3353 & tmp3357);
  wire tmp3359;
  assign tmp3359 = (tmp3332 & tmp3345) | (tmp3332 & tmp3358) | (tmp3345 & tmp3358);
  wire tmp3360;
  assign tmp3360 = 1'b0;
  wire tmp3361;
  assign tmp3361 = 1'b0;
  wire tmp3362;
  assign tmp3362 = 1'b0;
  wire tmp3363;
  assign tmp3363 = (tmp3360 & tmp3361) | (tmp3360 & tmp3362) | (tmp3361 & tmp3362);
  wire tmp3364;
  assign tmp3364 = 1'b0;
  wire tmp3365;
  assign tmp3365 = 1'b0;
  wire tmp3366;
  assign tmp3366 = 1'b0;
  wire tmp3367;
  assign tmp3367 = (tmp3364 & tmp3365) | (tmp3364 & tmp3366) | (tmp3365 & tmp3366);
  wire tmp3368;
  assign tmp3368 = 1'b0;
  wire tmp3369;
  assign tmp3369 = 1'b0;
  wire tmp3370;
  assign tmp3370 = 1'b0;
  wire tmp3371;
  assign tmp3371 = (tmp3368 & tmp3369) | (tmp3368 & tmp3370) | (tmp3369 & tmp3370);
  wire tmp3372;
  assign tmp3372 = (tmp3363 & tmp3367) | (tmp3363 & tmp3371) | (tmp3367 & tmp3371);
  wire tmp3373;
  assign tmp3373 = 1'b0;
  wire tmp3374;
  assign tmp3374 = 1'b0;
  wire tmp3375;
  assign tmp3375 = 1'b0;
  wire tmp3376;
  assign tmp3376 = (tmp3373 & tmp3374) | (tmp3373 & tmp3375) | (tmp3374 & tmp3375);
  wire tmp3377;
  assign tmp3377 = 1'b0;
  wire tmp3378;
  assign tmp3378 = 1'b1;
  wire tmp3379;
  assign tmp3379 = 1'b0;
  wire tmp3380;
  assign tmp3380 = (tmp3377 & tmp3378) | (tmp3377 & tmp3379) | (tmp3378 & tmp3379);
  wire tmp3381;
  assign tmp3381 = 1'b0;
  wire tmp3382;
  assign tmp3382 = 1'b0;
  wire tmp3383;
  assign tmp3383 = 1'b0;
  wire tmp3384;
  assign tmp3384 = (tmp3381 & tmp3382) | (tmp3381 & tmp3383) | (tmp3382 & tmp3383);
  wire tmp3385;
  assign tmp3385 = (tmp3376 & tmp3380) | (tmp3376 & tmp3384) | (tmp3380 & tmp3384);
  wire tmp3386;
  assign tmp3386 = 1'b0;
  wire tmp3387;
  assign tmp3387 = 1'b0;
  wire tmp3388;
  assign tmp3388 = 1'b0;
  wire tmp3389;
  assign tmp3389 = (tmp3386 & tmp3387) | (tmp3386 & tmp3388) | (tmp3387 & tmp3388);
  wire tmp3390;
  assign tmp3390 = 1'b0;
  wire tmp3391;
  assign tmp3391 = 1'b0;
  wire tmp3392;
  assign tmp3392 = 1'b0;
  wire tmp3393;
  assign tmp3393 = (tmp3390 & tmp3391) | (tmp3390 & tmp3392) | (tmp3391 & tmp3392);
  wire tmp3394;
  assign tmp3394 = 1'b0;
  wire tmp3395;
  assign tmp3395 = 1'b0;
  wire tmp3396;
  assign tmp3396 = 1'b0;
  wire tmp3397;
  assign tmp3397 = (tmp3394 & tmp3395) | (tmp3394 & tmp3396) | (tmp3395 & tmp3396);
  wire tmp3398;
  assign tmp3398 = (tmp3389 & tmp3393) | (tmp3389 & tmp3397) | (tmp3393 & tmp3397);
  wire tmp3399;
  assign tmp3399 = (tmp3372 & tmp3385) | (tmp3372 & tmp3398) | (tmp3385 & tmp3398);
  wire tmp3400;
  assign tmp3400 = (tmp3319 & tmp3359) | (tmp3319 & tmp3399) | (tmp3359 & tmp3399);
  wire tmp3401;
  assign tmp3401 = pi2;
  wire tmp3402;
  assign tmp3402 = pi3;
  wire tmp3403;
  assign tmp3403 = 1'b0;
  wire tmp3404;
  assign tmp3404 = (tmp3401 & tmp3402) | (tmp3401 & tmp3403) | (tmp3402 & tmp3403);
  wire tmp3405;
  assign tmp3405 = pi3;
  wire tmp3406;
  assign tmp3406 = 1'b1;
  wire tmp3407;
  assign tmp3407 = 1'b0;
  wire tmp3408;
  assign tmp3408 = (tmp3405 & tmp3406) | (tmp3405 & tmp3407) | (tmp3406 & tmp3407);
  wire tmp3409;
  assign tmp3409 = 1'b0;
  wire tmp3410;
  assign tmp3410 = 1'b0;
  wire tmp3411;
  assign tmp3411 = 1'b0;
  wire tmp3412;
  assign tmp3412 = (tmp3409 & tmp3410) | (tmp3409 & tmp3411) | (tmp3410 & tmp3411);
  wire tmp3413;
  assign tmp3413 = (tmp3404 & tmp3408) | (tmp3404 & tmp3412) | (tmp3408 & tmp3412);
  wire tmp3414;
  assign tmp3414 = pi3;
  wire tmp3415;
  assign tmp3415 = 1'b1;
  wire tmp3416;
  assign tmp3416 = 1'b0;
  wire tmp3417;
  assign tmp3417 = (tmp3414 & tmp3415) | (tmp3414 & tmp3416) | (tmp3415 & tmp3416);
  wire tmp3418;
  assign tmp3418 = 1'b1;
  wire tmp3419;
  assign tmp3419 = 1'b1;
  wire tmp3420;
  assign tmp3420 = 1'b1;
  wire tmp3421;
  assign tmp3421 = (tmp3418 & tmp3419) | (tmp3418 & tmp3420) | (tmp3419 & tmp3420);
  wire tmp3422;
  assign tmp3422 = 1'b0;
  wire tmp3423;
  assign tmp3423 = 1'b1;
  wire tmp3424;
  assign tmp3424 = 1'b0;
  wire tmp3425;
  assign tmp3425 = (tmp3422 & tmp3423) | (tmp3422 & tmp3424) | (tmp3423 & tmp3424);
  wire tmp3426;
  assign tmp3426 = (tmp3417 & tmp3421) | (tmp3417 & tmp3425) | (tmp3421 & tmp3425);
  wire tmp3427;
  assign tmp3427 = 1'b0;
  wire tmp3428;
  assign tmp3428 = 1'b0;
  wire tmp3429;
  assign tmp3429 = 1'b0;
  wire tmp3430;
  assign tmp3430 = (tmp3427 & tmp3428) | (tmp3427 & tmp3429) | (tmp3428 & tmp3429);
  wire tmp3431;
  assign tmp3431 = 1'b0;
  wire tmp3432;
  assign tmp3432 = 1'b1;
  wire tmp3433;
  assign tmp3433 = 1'b0;
  wire tmp3434;
  assign tmp3434 = (tmp3431 & tmp3432) | (tmp3431 & tmp3433) | (tmp3432 & tmp3433);
  wire tmp3435;
  assign tmp3435 = 1'b0;
  wire tmp3436;
  assign tmp3436 = 1'b0;
  wire tmp3437;
  assign tmp3437 = 1'b0;
  wire tmp3438;
  assign tmp3438 = (tmp3435 & tmp3436) | (tmp3435 & tmp3437) | (tmp3436 & tmp3437);
  wire tmp3439;
  assign tmp3439 = (tmp3430 & tmp3434) | (tmp3430 & tmp3438) | (tmp3434 & tmp3438);
  wire tmp3440;
  assign tmp3440 = (tmp3413 & tmp3426) | (tmp3413 & tmp3439) | (tmp3426 & tmp3439);
  wire tmp3441;
  assign tmp3441 = pi3;
  wire tmp3442;
  assign tmp3442 = 1'b1;
  wire tmp3443;
  assign tmp3443 = 1'b0;
  wire tmp3444;
  assign tmp3444 = (tmp3441 & tmp3442) | (tmp3441 & tmp3443) | (tmp3442 & tmp3443);
  wire tmp3445;
  assign tmp3445 = 1'b1;
  wire tmp3446;
  assign tmp3446 = 1'b1;
  wire tmp3447;
  assign tmp3447 = 1'b1;
  wire tmp3448;
  assign tmp3448 = (tmp3445 & tmp3446) | (tmp3445 & tmp3447) | (tmp3446 & tmp3447);
  wire tmp3449;
  assign tmp3449 = 1'b0;
  wire tmp3450;
  assign tmp3450 = 1'b1;
  wire tmp3451;
  assign tmp3451 = 1'b0;
  wire tmp3452;
  assign tmp3452 = (tmp3449 & tmp3450) | (tmp3449 & tmp3451) | (tmp3450 & tmp3451);
  wire tmp3453;
  assign tmp3453 = (tmp3444 & tmp3448) | (tmp3444 & tmp3452) | (tmp3448 & tmp3452);
  wire tmp3454;
  assign tmp3454 = 1'b1;
  wire tmp3455;
  assign tmp3455 = 1'b1;
  wire tmp3456;
  assign tmp3456 = 1'b1;
  wire tmp3457;
  assign tmp3457 = (tmp3454 & tmp3455) | (tmp3454 & tmp3456) | (tmp3455 & tmp3456);
  wire tmp3458;
  assign tmp3458 = 1'b1;
  wire tmp3459;
  assign tmp3459 = 1'b1;
  wire tmp3460;
  assign tmp3460 = 1'b1;
  wire tmp3461;
  assign tmp3461 = (tmp3458 & tmp3459) | (tmp3458 & tmp3460) | (tmp3459 & tmp3460);
  wire tmp3462;
  assign tmp3462 = 1'b1;
  wire tmp3463;
  assign tmp3463 = 1'b1;
  wire tmp3464;
  assign tmp3464 = 1'b1;
  wire tmp3465;
  assign tmp3465 = (tmp3462 & tmp3463) | (tmp3462 & tmp3464) | (tmp3463 & tmp3464);
  wire tmp3466;
  assign tmp3466 = (tmp3457 & tmp3461) | (tmp3457 & tmp3465) | (tmp3461 & tmp3465);
  wire tmp3467;
  assign tmp3467 = 1'b0;
  wire tmp3468;
  assign tmp3468 = 1'b1;
  wire tmp3469;
  assign tmp3469 = 1'b0;
  wire tmp3470;
  assign tmp3470 = (tmp3467 & tmp3468) | (tmp3467 & tmp3469) | (tmp3468 & tmp3469);
  wire tmp3471;
  assign tmp3471 = 1'b1;
  wire tmp3472;
  assign tmp3472 = 1'b1;
  wire tmp3473;
  assign tmp3473 = 1'b1;
  wire tmp3474;
  assign tmp3474 = (tmp3471 & tmp3472) | (tmp3471 & tmp3473) | (tmp3472 & tmp3473);
  wire tmp3475;
  assign tmp3475 = 1'b0;
  wire tmp3476;
  assign tmp3476 = 1'b1;
  wire tmp3477;
  assign tmp3477 = 1'b0;
  wire tmp3478;
  assign tmp3478 = (tmp3475 & tmp3476) | (tmp3475 & tmp3477) | (tmp3476 & tmp3477);
  wire tmp3479;
  assign tmp3479 = (tmp3470 & tmp3474) | (tmp3470 & tmp3478) | (tmp3474 & tmp3478);
  wire tmp3480;
  assign tmp3480 = (tmp3453 & tmp3466) | (tmp3453 & tmp3479) | (tmp3466 & tmp3479);
  wire tmp3481;
  assign tmp3481 = 1'b0;
  wire tmp3482;
  assign tmp3482 = 1'b0;
  wire tmp3483;
  assign tmp3483 = 1'b0;
  wire tmp3484;
  assign tmp3484 = (tmp3481 & tmp3482) | (tmp3481 & tmp3483) | (tmp3482 & tmp3483);
  wire tmp3485;
  assign tmp3485 = 1'b0;
  wire tmp3486;
  assign tmp3486 = 1'b1;
  wire tmp3487;
  assign tmp3487 = 1'b0;
  wire tmp3488;
  assign tmp3488 = (tmp3485 & tmp3486) | (tmp3485 & tmp3487) | (tmp3486 & tmp3487);
  wire tmp3489;
  assign tmp3489 = 1'b0;
  wire tmp3490;
  assign tmp3490 = 1'b0;
  wire tmp3491;
  assign tmp3491 = 1'b0;
  wire tmp3492;
  assign tmp3492 = (tmp3489 & tmp3490) | (tmp3489 & tmp3491) | (tmp3490 & tmp3491);
  wire tmp3493;
  assign tmp3493 = (tmp3484 & tmp3488) | (tmp3484 & tmp3492) | (tmp3488 & tmp3492);
  wire tmp3494;
  assign tmp3494 = 1'b0;
  wire tmp3495;
  assign tmp3495 = 1'b1;
  wire tmp3496;
  assign tmp3496 = 1'b0;
  wire tmp3497;
  assign tmp3497 = (tmp3494 & tmp3495) | (tmp3494 & tmp3496) | (tmp3495 & tmp3496);
  wire tmp3498;
  assign tmp3498 = 1'b1;
  wire tmp3499;
  assign tmp3499 = 1'b1;
  wire tmp3500;
  assign tmp3500 = 1'b1;
  wire tmp3501;
  assign tmp3501 = (tmp3498 & tmp3499) | (tmp3498 & tmp3500) | (tmp3499 & tmp3500);
  wire tmp3502;
  assign tmp3502 = 1'b0;
  wire tmp3503;
  assign tmp3503 = 1'b1;
  wire tmp3504;
  assign tmp3504 = 1'b0;
  wire tmp3505;
  assign tmp3505 = (tmp3502 & tmp3503) | (tmp3502 & tmp3504) | (tmp3503 & tmp3504);
  wire tmp3506;
  assign tmp3506 = (tmp3497 & tmp3501) | (tmp3497 & tmp3505) | (tmp3501 & tmp3505);
  wire tmp3507;
  assign tmp3507 = 1'b0;
  wire tmp3508;
  assign tmp3508 = 1'b0;
  wire tmp3509;
  assign tmp3509 = 1'b0;
  wire tmp3510;
  assign tmp3510 = (tmp3507 & tmp3508) | (tmp3507 & tmp3509) | (tmp3508 & tmp3509);
  wire tmp3511;
  assign tmp3511 = 1'b0;
  wire tmp3512;
  assign tmp3512 = 1'b1;
  wire tmp3513;
  assign tmp3513 = 1'b0;
  wire tmp3514;
  assign tmp3514 = (tmp3511 & tmp3512) | (tmp3511 & tmp3513) | (tmp3512 & tmp3513);
  wire tmp3515;
  assign tmp3515 = 1'b0;
  wire tmp3516;
  assign tmp3516 = 1'b0;
  wire tmp3517;
  assign tmp3517 = 1'b0;
  wire tmp3518;
  assign tmp3518 = (tmp3515 & tmp3516) | (tmp3515 & tmp3517) | (tmp3516 & tmp3517);
  wire tmp3519;
  assign tmp3519 = (tmp3510 & tmp3514) | (tmp3510 & tmp3518) | (tmp3514 & tmp3518);
  wire tmp3520;
  assign tmp3520 = (tmp3493 & tmp3506) | (tmp3493 & tmp3519) | (tmp3506 & tmp3519);
  wire tmp3521;
  assign tmp3521 = (tmp3440 & tmp3480) | (tmp3440 & tmp3520) | (tmp3480 & tmp3520);
  wire tmp3522;
  assign tmp3522 = 1'b0;
  wire tmp3523;
  assign tmp3523 = 1'b0;
  wire tmp3524;
  assign tmp3524 = 1'b0;
  wire tmp3525;
  assign tmp3525 = (tmp3522 & tmp3523) | (tmp3522 & tmp3524) | (tmp3523 & tmp3524);
  wire tmp3526;
  assign tmp3526 = 1'b0;
  wire tmp3527;
  assign tmp3527 = 1'b0;
  wire tmp3528;
  assign tmp3528 = 1'b0;
  wire tmp3529;
  assign tmp3529 = (tmp3526 & tmp3527) | (tmp3526 & tmp3528) | (tmp3527 & tmp3528);
  wire tmp3530;
  assign tmp3530 = 1'b0;
  wire tmp3531;
  assign tmp3531 = 1'b0;
  wire tmp3532;
  assign tmp3532 = 1'b0;
  wire tmp3533;
  assign tmp3533 = (tmp3530 & tmp3531) | (tmp3530 & tmp3532) | (tmp3531 & tmp3532);
  wire tmp3534;
  assign tmp3534 = (tmp3525 & tmp3529) | (tmp3525 & tmp3533) | (tmp3529 & tmp3533);
  wire tmp3535;
  assign tmp3535 = 1'b0;
  wire tmp3536;
  assign tmp3536 = 1'b0;
  wire tmp3537;
  assign tmp3537 = 1'b0;
  wire tmp3538;
  assign tmp3538 = (tmp3535 & tmp3536) | (tmp3535 & tmp3537) | (tmp3536 & tmp3537);
  wire tmp3539;
  assign tmp3539 = 1'b0;
  wire tmp3540;
  assign tmp3540 = 1'b1;
  wire tmp3541;
  assign tmp3541 = 1'b0;
  wire tmp3542;
  assign tmp3542 = (tmp3539 & tmp3540) | (tmp3539 & tmp3541) | (tmp3540 & tmp3541);
  wire tmp3543;
  assign tmp3543 = 1'b0;
  wire tmp3544;
  assign tmp3544 = 1'b0;
  wire tmp3545;
  assign tmp3545 = 1'b0;
  wire tmp3546;
  assign tmp3546 = (tmp3543 & tmp3544) | (tmp3543 & tmp3545) | (tmp3544 & tmp3545);
  wire tmp3547;
  assign tmp3547 = (tmp3538 & tmp3542) | (tmp3538 & tmp3546) | (tmp3542 & tmp3546);
  wire tmp3548;
  assign tmp3548 = 1'b0;
  wire tmp3549;
  assign tmp3549 = 1'b0;
  wire tmp3550;
  assign tmp3550 = 1'b0;
  wire tmp3551;
  assign tmp3551 = (tmp3548 & tmp3549) | (tmp3548 & tmp3550) | (tmp3549 & tmp3550);
  wire tmp3552;
  assign tmp3552 = 1'b0;
  wire tmp3553;
  assign tmp3553 = 1'b0;
  wire tmp3554;
  assign tmp3554 = 1'b0;
  wire tmp3555;
  assign tmp3555 = (tmp3552 & tmp3553) | (tmp3552 & tmp3554) | (tmp3553 & tmp3554);
  wire tmp3556;
  assign tmp3556 = 1'b0;
  wire tmp3557;
  assign tmp3557 = 1'b0;
  wire tmp3558;
  assign tmp3558 = 1'b0;
  wire tmp3559;
  assign tmp3559 = (tmp3556 & tmp3557) | (tmp3556 & tmp3558) | (tmp3557 & tmp3558);
  wire tmp3560;
  assign tmp3560 = (tmp3551 & tmp3555) | (tmp3551 & tmp3559) | (tmp3555 & tmp3559);
  wire tmp3561;
  assign tmp3561 = (tmp3534 & tmp3547) | (tmp3534 & tmp3560) | (tmp3547 & tmp3560);
  wire tmp3562;
  assign tmp3562 = 1'b0;
  wire tmp3563;
  assign tmp3563 = 1'b0;
  wire tmp3564;
  assign tmp3564 = 1'b0;
  wire tmp3565;
  assign tmp3565 = (tmp3562 & tmp3563) | (tmp3562 & tmp3564) | (tmp3563 & tmp3564);
  wire tmp3566;
  assign tmp3566 = 1'b0;
  wire tmp3567;
  assign tmp3567 = 1'b1;
  wire tmp3568;
  assign tmp3568 = 1'b0;
  wire tmp3569;
  assign tmp3569 = (tmp3566 & tmp3567) | (tmp3566 & tmp3568) | (tmp3567 & tmp3568);
  wire tmp3570;
  assign tmp3570 = 1'b0;
  wire tmp3571;
  assign tmp3571 = 1'b0;
  wire tmp3572;
  assign tmp3572 = 1'b0;
  wire tmp3573;
  assign tmp3573 = (tmp3570 & tmp3571) | (tmp3570 & tmp3572) | (tmp3571 & tmp3572);
  wire tmp3574;
  assign tmp3574 = (tmp3565 & tmp3569) | (tmp3565 & tmp3573) | (tmp3569 & tmp3573);
  wire tmp3575;
  assign tmp3575 = 1'b0;
  wire tmp3576;
  assign tmp3576 = 1'b1;
  wire tmp3577;
  assign tmp3577 = 1'b0;
  wire tmp3578;
  assign tmp3578 = (tmp3575 & tmp3576) | (tmp3575 & tmp3577) | (tmp3576 & tmp3577);
  wire tmp3579;
  assign tmp3579 = 1'b1;
  wire tmp3580;
  assign tmp3580 = 1'b1;
  wire tmp3581;
  assign tmp3581 = 1'b1;
  wire tmp3582;
  assign tmp3582 = (tmp3579 & tmp3580) | (tmp3579 & tmp3581) | (tmp3580 & tmp3581);
  wire tmp3583;
  assign tmp3583 = 1'b0;
  wire tmp3584;
  assign tmp3584 = 1'b1;
  wire tmp3585;
  assign tmp3585 = 1'b0;
  wire tmp3586;
  assign tmp3586 = (tmp3583 & tmp3584) | (tmp3583 & tmp3585) | (tmp3584 & tmp3585);
  wire tmp3587;
  assign tmp3587 = (tmp3578 & tmp3582) | (tmp3578 & tmp3586) | (tmp3582 & tmp3586);
  wire tmp3588;
  assign tmp3588 = 1'b0;
  wire tmp3589;
  assign tmp3589 = 1'b0;
  wire tmp3590;
  assign tmp3590 = 1'b0;
  wire tmp3591;
  assign tmp3591 = (tmp3588 & tmp3589) | (tmp3588 & tmp3590) | (tmp3589 & tmp3590);
  wire tmp3592;
  assign tmp3592 = 1'b0;
  wire tmp3593;
  assign tmp3593 = 1'b1;
  wire tmp3594;
  assign tmp3594 = 1'b0;
  wire tmp3595;
  assign tmp3595 = (tmp3592 & tmp3593) | (tmp3592 & tmp3594) | (tmp3593 & tmp3594);
  wire tmp3596;
  assign tmp3596 = 1'b0;
  wire tmp3597;
  assign tmp3597 = 1'b0;
  wire tmp3598;
  assign tmp3598 = 1'b0;
  wire tmp3599;
  assign tmp3599 = (tmp3596 & tmp3597) | (tmp3596 & tmp3598) | (tmp3597 & tmp3598);
  wire tmp3600;
  assign tmp3600 = (tmp3591 & tmp3595) | (tmp3591 & tmp3599) | (tmp3595 & tmp3599);
  wire tmp3601;
  assign tmp3601 = (tmp3574 & tmp3587) | (tmp3574 & tmp3600) | (tmp3587 & tmp3600);
  wire tmp3602;
  assign tmp3602 = 1'b0;
  wire tmp3603;
  assign tmp3603 = 1'b0;
  wire tmp3604;
  assign tmp3604 = 1'b0;
  wire tmp3605;
  assign tmp3605 = (tmp3602 & tmp3603) | (tmp3602 & tmp3604) | (tmp3603 & tmp3604);
  wire tmp3606;
  assign tmp3606 = 1'b0;
  wire tmp3607;
  assign tmp3607 = 1'b0;
  wire tmp3608;
  assign tmp3608 = 1'b0;
  wire tmp3609;
  assign tmp3609 = (tmp3606 & tmp3607) | (tmp3606 & tmp3608) | (tmp3607 & tmp3608);
  wire tmp3610;
  assign tmp3610 = 1'b0;
  wire tmp3611;
  assign tmp3611 = 1'b0;
  wire tmp3612;
  assign tmp3612 = 1'b0;
  wire tmp3613;
  assign tmp3613 = (tmp3610 & tmp3611) | (tmp3610 & tmp3612) | (tmp3611 & tmp3612);
  wire tmp3614;
  assign tmp3614 = (tmp3605 & tmp3609) | (tmp3605 & tmp3613) | (tmp3609 & tmp3613);
  wire tmp3615;
  assign tmp3615 = 1'b0;
  wire tmp3616;
  assign tmp3616 = 1'b0;
  wire tmp3617;
  assign tmp3617 = 1'b0;
  wire tmp3618;
  assign tmp3618 = (tmp3615 & tmp3616) | (tmp3615 & tmp3617) | (tmp3616 & tmp3617);
  wire tmp3619;
  assign tmp3619 = 1'b0;
  wire tmp3620;
  assign tmp3620 = 1'b1;
  wire tmp3621;
  assign tmp3621 = 1'b0;
  wire tmp3622;
  assign tmp3622 = (tmp3619 & tmp3620) | (tmp3619 & tmp3621) | (tmp3620 & tmp3621);
  wire tmp3623;
  assign tmp3623 = 1'b0;
  wire tmp3624;
  assign tmp3624 = 1'b0;
  wire tmp3625;
  assign tmp3625 = 1'b0;
  wire tmp3626;
  assign tmp3626 = (tmp3623 & tmp3624) | (tmp3623 & tmp3625) | (tmp3624 & tmp3625);
  wire tmp3627;
  assign tmp3627 = (tmp3618 & tmp3622) | (tmp3618 & tmp3626) | (tmp3622 & tmp3626);
  wire tmp3628;
  assign tmp3628 = 1'b0;
  wire tmp3629;
  assign tmp3629 = 1'b0;
  wire tmp3630;
  assign tmp3630 = 1'b0;
  wire tmp3631;
  assign tmp3631 = (tmp3628 & tmp3629) | (tmp3628 & tmp3630) | (tmp3629 & tmp3630);
  wire tmp3632;
  assign tmp3632 = 1'b0;
  wire tmp3633;
  assign tmp3633 = 1'b0;
  wire tmp3634;
  assign tmp3634 = 1'b0;
  wire tmp3635;
  assign tmp3635 = (tmp3632 & tmp3633) | (tmp3632 & tmp3634) | (tmp3633 & tmp3634);
  wire tmp3636;
  assign tmp3636 = 1'b0;
  wire tmp3637;
  assign tmp3637 = 1'b0;
  wire tmp3638;
  assign tmp3638 = 1'b0;
  wire tmp3639;
  assign tmp3639 = (tmp3636 & tmp3637) | (tmp3636 & tmp3638) | (tmp3637 & tmp3638);
  wire tmp3640;
  assign tmp3640 = (tmp3631 & tmp3635) | (tmp3631 & tmp3639) | (tmp3635 & tmp3639);
  wire tmp3641;
  assign tmp3641 = (tmp3614 & tmp3627) | (tmp3614 & tmp3640) | (tmp3627 & tmp3640);
  wire tmp3642;
  assign tmp3642 = (tmp3561 & tmp3601) | (tmp3561 & tmp3641) | (tmp3601 & tmp3641);
  wire tmp3643;
  assign tmp3643 = (tmp3400 & tmp3521) | (tmp3400 & tmp3642) | (tmp3521 & tmp3642);
  wire tmp3644;
  assign tmp3644 = pi2;
  wire tmp3645;
  assign tmp3645 = pi3;
  wire tmp3646;
  assign tmp3646 = 1'b0;
  wire tmp3647;
  assign tmp3647 = (tmp3644 & tmp3645) | (tmp3644 & tmp3646) | (tmp3645 & tmp3646);
  wire tmp3648;
  assign tmp3648 = pi3;
  wire tmp3649;
  assign tmp3649 = 1'b1;
  wire tmp3650;
  assign tmp3650 = 1'b0;
  wire tmp3651;
  assign tmp3651 = (tmp3648 & tmp3649) | (tmp3648 & tmp3650) | (tmp3649 & tmp3650);
  wire tmp3652;
  assign tmp3652 = 1'b0;
  wire tmp3653;
  assign tmp3653 = 1'b0;
  wire tmp3654;
  assign tmp3654 = 1'b0;
  wire tmp3655;
  assign tmp3655 = (tmp3652 & tmp3653) | (tmp3652 & tmp3654) | (tmp3653 & tmp3654);
  wire tmp3656;
  assign tmp3656 = (tmp3647 & tmp3651) | (tmp3647 & tmp3655) | (tmp3651 & tmp3655);
  wire tmp3657;
  assign tmp3657 = pi3;
  wire tmp3658;
  assign tmp3658 = 1'b1;
  wire tmp3659;
  assign tmp3659 = 1'b0;
  wire tmp3660;
  assign tmp3660 = (tmp3657 & tmp3658) | (tmp3657 & tmp3659) | (tmp3658 & tmp3659);
  wire tmp3661;
  assign tmp3661 = 1'b1;
  wire tmp3662;
  assign tmp3662 = 1'b1;
  wire tmp3663;
  assign tmp3663 = 1'b1;
  wire tmp3664;
  assign tmp3664 = (tmp3661 & tmp3662) | (tmp3661 & tmp3663) | (tmp3662 & tmp3663);
  wire tmp3665;
  assign tmp3665 = 1'b0;
  wire tmp3666;
  assign tmp3666 = 1'b1;
  wire tmp3667;
  assign tmp3667 = 1'b0;
  wire tmp3668;
  assign tmp3668 = (tmp3665 & tmp3666) | (tmp3665 & tmp3667) | (tmp3666 & tmp3667);
  wire tmp3669;
  assign tmp3669 = (tmp3660 & tmp3664) | (tmp3660 & tmp3668) | (tmp3664 & tmp3668);
  wire tmp3670;
  assign tmp3670 = 1'b0;
  wire tmp3671;
  assign tmp3671 = 1'b0;
  wire tmp3672;
  assign tmp3672 = 1'b0;
  wire tmp3673;
  assign tmp3673 = (tmp3670 & tmp3671) | (tmp3670 & tmp3672) | (tmp3671 & tmp3672);
  wire tmp3674;
  assign tmp3674 = 1'b0;
  wire tmp3675;
  assign tmp3675 = 1'b1;
  wire tmp3676;
  assign tmp3676 = 1'b0;
  wire tmp3677;
  assign tmp3677 = (tmp3674 & tmp3675) | (tmp3674 & tmp3676) | (tmp3675 & tmp3676);
  wire tmp3678;
  assign tmp3678 = 1'b0;
  wire tmp3679;
  assign tmp3679 = 1'b0;
  wire tmp3680;
  assign tmp3680 = 1'b0;
  wire tmp3681;
  assign tmp3681 = (tmp3678 & tmp3679) | (tmp3678 & tmp3680) | (tmp3679 & tmp3680);
  wire tmp3682;
  assign tmp3682 = (tmp3673 & tmp3677) | (tmp3673 & tmp3681) | (tmp3677 & tmp3681);
  wire tmp3683;
  assign tmp3683 = (tmp3656 & tmp3669) | (tmp3656 & tmp3682) | (tmp3669 & tmp3682);
  wire tmp3684;
  assign tmp3684 = pi3;
  wire tmp3685;
  assign tmp3685 = 1'b1;
  wire tmp3686;
  assign tmp3686 = 1'b0;
  wire tmp3687;
  assign tmp3687 = (tmp3684 & tmp3685) | (tmp3684 & tmp3686) | (tmp3685 & tmp3686);
  wire tmp3688;
  assign tmp3688 = 1'b1;
  wire tmp3689;
  assign tmp3689 = 1'b1;
  wire tmp3690;
  assign tmp3690 = 1'b1;
  wire tmp3691;
  assign tmp3691 = (tmp3688 & tmp3689) | (tmp3688 & tmp3690) | (tmp3689 & tmp3690);
  wire tmp3692;
  assign tmp3692 = 1'b0;
  wire tmp3693;
  assign tmp3693 = 1'b1;
  wire tmp3694;
  assign tmp3694 = 1'b0;
  wire tmp3695;
  assign tmp3695 = (tmp3692 & tmp3693) | (tmp3692 & tmp3694) | (tmp3693 & tmp3694);
  wire tmp3696;
  assign tmp3696 = (tmp3687 & tmp3691) | (tmp3687 & tmp3695) | (tmp3691 & tmp3695);
  wire tmp3697;
  assign tmp3697 = 1'b1;
  wire tmp3698;
  assign tmp3698 = 1'b1;
  wire tmp3699;
  assign tmp3699 = 1'b1;
  wire tmp3700;
  assign tmp3700 = (tmp3697 & tmp3698) | (tmp3697 & tmp3699) | (tmp3698 & tmp3699);
  wire tmp3701;
  assign tmp3701 = 1'b1;
  wire tmp3702;
  assign tmp3702 = 1'b1;
  wire tmp3703;
  assign tmp3703 = 1'b1;
  wire tmp3704;
  assign tmp3704 = (tmp3701 & tmp3702) | (tmp3701 & tmp3703) | (tmp3702 & tmp3703);
  wire tmp3705;
  assign tmp3705 = 1'b1;
  wire tmp3706;
  assign tmp3706 = 1'b1;
  wire tmp3707;
  assign tmp3707 = 1'b1;
  wire tmp3708;
  assign tmp3708 = (tmp3705 & tmp3706) | (tmp3705 & tmp3707) | (tmp3706 & tmp3707);
  wire tmp3709;
  assign tmp3709 = (tmp3700 & tmp3704) | (tmp3700 & tmp3708) | (tmp3704 & tmp3708);
  wire tmp3710;
  assign tmp3710 = 1'b0;
  wire tmp3711;
  assign tmp3711 = 1'b1;
  wire tmp3712;
  assign tmp3712 = 1'b0;
  wire tmp3713;
  assign tmp3713 = (tmp3710 & tmp3711) | (tmp3710 & tmp3712) | (tmp3711 & tmp3712);
  wire tmp3714;
  assign tmp3714 = 1'b1;
  wire tmp3715;
  assign tmp3715 = 1'b1;
  wire tmp3716;
  assign tmp3716 = 1'b1;
  wire tmp3717;
  assign tmp3717 = (tmp3714 & tmp3715) | (tmp3714 & tmp3716) | (tmp3715 & tmp3716);
  wire tmp3718;
  assign tmp3718 = 1'b0;
  wire tmp3719;
  assign tmp3719 = 1'b1;
  wire tmp3720;
  assign tmp3720 = 1'b0;
  wire tmp3721;
  assign tmp3721 = (tmp3718 & tmp3719) | (tmp3718 & tmp3720) | (tmp3719 & tmp3720);
  wire tmp3722;
  assign tmp3722 = (tmp3713 & tmp3717) | (tmp3713 & tmp3721) | (tmp3717 & tmp3721);
  wire tmp3723;
  assign tmp3723 = (tmp3696 & tmp3709) | (tmp3696 & tmp3722) | (tmp3709 & tmp3722);
  wire tmp3724;
  assign tmp3724 = 1'b0;
  wire tmp3725;
  assign tmp3725 = 1'b0;
  wire tmp3726;
  assign tmp3726 = 1'b0;
  wire tmp3727;
  assign tmp3727 = (tmp3724 & tmp3725) | (tmp3724 & tmp3726) | (tmp3725 & tmp3726);
  wire tmp3728;
  assign tmp3728 = 1'b0;
  wire tmp3729;
  assign tmp3729 = 1'b1;
  wire tmp3730;
  assign tmp3730 = 1'b0;
  wire tmp3731;
  assign tmp3731 = (tmp3728 & tmp3729) | (tmp3728 & tmp3730) | (tmp3729 & tmp3730);
  wire tmp3732;
  assign tmp3732 = 1'b0;
  wire tmp3733;
  assign tmp3733 = 1'b0;
  wire tmp3734;
  assign tmp3734 = 1'b0;
  wire tmp3735;
  assign tmp3735 = (tmp3732 & tmp3733) | (tmp3732 & tmp3734) | (tmp3733 & tmp3734);
  wire tmp3736;
  assign tmp3736 = (tmp3727 & tmp3731) | (tmp3727 & tmp3735) | (tmp3731 & tmp3735);
  wire tmp3737;
  assign tmp3737 = 1'b0;
  wire tmp3738;
  assign tmp3738 = 1'b1;
  wire tmp3739;
  assign tmp3739 = 1'b0;
  wire tmp3740;
  assign tmp3740 = (tmp3737 & tmp3738) | (tmp3737 & tmp3739) | (tmp3738 & tmp3739);
  wire tmp3741;
  assign tmp3741 = 1'b1;
  wire tmp3742;
  assign tmp3742 = 1'b1;
  wire tmp3743;
  assign tmp3743 = 1'b1;
  wire tmp3744;
  assign tmp3744 = (tmp3741 & tmp3742) | (tmp3741 & tmp3743) | (tmp3742 & tmp3743);
  wire tmp3745;
  assign tmp3745 = 1'b0;
  wire tmp3746;
  assign tmp3746 = 1'b1;
  wire tmp3747;
  assign tmp3747 = 1'b0;
  wire tmp3748;
  assign tmp3748 = (tmp3745 & tmp3746) | (tmp3745 & tmp3747) | (tmp3746 & tmp3747);
  wire tmp3749;
  assign tmp3749 = (tmp3740 & tmp3744) | (tmp3740 & tmp3748) | (tmp3744 & tmp3748);
  wire tmp3750;
  assign tmp3750 = 1'b0;
  wire tmp3751;
  assign tmp3751 = 1'b0;
  wire tmp3752;
  assign tmp3752 = 1'b0;
  wire tmp3753;
  assign tmp3753 = (tmp3750 & tmp3751) | (tmp3750 & tmp3752) | (tmp3751 & tmp3752);
  wire tmp3754;
  assign tmp3754 = 1'b0;
  wire tmp3755;
  assign tmp3755 = 1'b1;
  wire tmp3756;
  assign tmp3756 = 1'b0;
  wire tmp3757;
  assign tmp3757 = (tmp3754 & tmp3755) | (tmp3754 & tmp3756) | (tmp3755 & tmp3756);
  wire tmp3758;
  assign tmp3758 = 1'b0;
  wire tmp3759;
  assign tmp3759 = 1'b0;
  wire tmp3760;
  assign tmp3760 = 1'b0;
  wire tmp3761;
  assign tmp3761 = (tmp3758 & tmp3759) | (tmp3758 & tmp3760) | (tmp3759 & tmp3760);
  wire tmp3762;
  assign tmp3762 = (tmp3753 & tmp3757) | (tmp3753 & tmp3761) | (tmp3757 & tmp3761);
  wire tmp3763;
  assign tmp3763 = (tmp3736 & tmp3749) | (tmp3736 & tmp3762) | (tmp3749 & tmp3762);
  wire tmp3764;
  assign tmp3764 = (tmp3683 & tmp3723) | (tmp3683 & tmp3763) | (tmp3723 & tmp3763);
  wire tmp3765;
  assign tmp3765 = pi3;
  wire tmp3766;
  assign tmp3766 = 1'b1;
  wire tmp3767;
  assign tmp3767 = 1'b0;
  wire tmp3768;
  assign tmp3768 = (tmp3765 & tmp3766) | (tmp3765 & tmp3767) | (tmp3766 & tmp3767);
  wire tmp3769;
  assign tmp3769 = 1'b1;
  wire tmp3770;
  assign tmp3770 = 1'b1;
  wire tmp3771;
  assign tmp3771 = 1'b1;
  wire tmp3772;
  assign tmp3772 = (tmp3769 & tmp3770) | (tmp3769 & tmp3771) | (tmp3770 & tmp3771);
  wire tmp3773;
  assign tmp3773 = 1'b0;
  wire tmp3774;
  assign tmp3774 = 1'b1;
  wire tmp3775;
  assign tmp3775 = 1'b0;
  wire tmp3776;
  assign tmp3776 = (tmp3773 & tmp3774) | (tmp3773 & tmp3775) | (tmp3774 & tmp3775);
  wire tmp3777;
  assign tmp3777 = (tmp3768 & tmp3772) | (tmp3768 & tmp3776) | (tmp3772 & tmp3776);
  wire tmp3778;
  assign tmp3778 = 1'b1;
  wire tmp3779;
  assign tmp3779 = 1'b1;
  wire tmp3780;
  assign tmp3780 = 1'b1;
  wire tmp3781;
  assign tmp3781 = (tmp3778 & tmp3779) | (tmp3778 & tmp3780) | (tmp3779 & tmp3780);
  wire tmp3782;
  assign tmp3782 = 1'b1;
  wire tmp3783;
  assign tmp3783 = 1'b1;
  wire tmp3784;
  assign tmp3784 = 1'b1;
  wire tmp3785;
  assign tmp3785 = (tmp3782 & tmp3783) | (tmp3782 & tmp3784) | (tmp3783 & tmp3784);
  wire tmp3786;
  assign tmp3786 = 1'b1;
  wire tmp3787;
  assign tmp3787 = 1'b1;
  wire tmp3788;
  assign tmp3788 = 1'b1;
  wire tmp3789;
  assign tmp3789 = (tmp3786 & tmp3787) | (tmp3786 & tmp3788) | (tmp3787 & tmp3788);
  wire tmp3790;
  assign tmp3790 = (tmp3781 & tmp3785) | (tmp3781 & tmp3789) | (tmp3785 & tmp3789);
  wire tmp3791;
  assign tmp3791 = 1'b0;
  wire tmp3792;
  assign tmp3792 = 1'b1;
  wire tmp3793;
  assign tmp3793 = 1'b0;
  wire tmp3794;
  assign tmp3794 = (tmp3791 & tmp3792) | (tmp3791 & tmp3793) | (tmp3792 & tmp3793);
  wire tmp3795;
  assign tmp3795 = 1'b1;
  wire tmp3796;
  assign tmp3796 = 1'b1;
  wire tmp3797;
  assign tmp3797 = 1'b1;
  wire tmp3798;
  assign tmp3798 = (tmp3795 & tmp3796) | (tmp3795 & tmp3797) | (tmp3796 & tmp3797);
  wire tmp3799;
  assign tmp3799 = 1'b0;
  wire tmp3800;
  assign tmp3800 = 1'b1;
  wire tmp3801;
  assign tmp3801 = 1'b0;
  wire tmp3802;
  assign tmp3802 = (tmp3799 & tmp3800) | (tmp3799 & tmp3801) | (tmp3800 & tmp3801);
  wire tmp3803;
  assign tmp3803 = (tmp3794 & tmp3798) | (tmp3794 & tmp3802) | (tmp3798 & tmp3802);
  wire tmp3804;
  assign tmp3804 = (tmp3777 & tmp3790) | (tmp3777 & tmp3803) | (tmp3790 & tmp3803);
  wire tmp3805;
  assign tmp3805 = 1'b1;
  wire tmp3806;
  assign tmp3806 = 1'b1;
  wire tmp3807;
  assign tmp3807 = 1'b1;
  wire tmp3808;
  assign tmp3808 = (tmp3805 & tmp3806) | (tmp3805 & tmp3807) | (tmp3806 & tmp3807);
  wire tmp3809;
  assign tmp3809 = 1'b1;
  wire tmp3810;
  assign tmp3810 = 1'b1;
  wire tmp3811;
  assign tmp3811 = 1'b1;
  wire tmp3812;
  assign tmp3812 = (tmp3809 & tmp3810) | (tmp3809 & tmp3811) | (tmp3810 & tmp3811);
  wire tmp3813;
  assign tmp3813 = 1'b1;
  wire tmp3814;
  assign tmp3814 = 1'b1;
  wire tmp3815;
  assign tmp3815 = 1'b1;
  wire tmp3816;
  assign tmp3816 = (tmp3813 & tmp3814) | (tmp3813 & tmp3815) | (tmp3814 & tmp3815);
  wire tmp3817;
  assign tmp3817 = (tmp3808 & tmp3812) | (tmp3808 & tmp3816) | (tmp3812 & tmp3816);
  wire tmp3818;
  assign tmp3818 = 1'b1;
  wire tmp3819;
  assign tmp3819 = 1'b1;
  wire tmp3820;
  assign tmp3820 = 1'b1;
  wire tmp3821;
  assign tmp3821 = (tmp3818 & tmp3819) | (tmp3818 & tmp3820) | (tmp3819 & tmp3820);
  wire tmp3822;
  assign tmp3822 = 1'b1;
  wire tmp3823;
  assign tmp3823 = ~pi4;
  wire tmp3824;
  assign tmp3824 = ~pi5;
  wire tmp3825;
  assign tmp3825 = (tmp3822 & tmp3823) | (tmp3822 & tmp3824) | (tmp3823 & tmp3824);
  wire tmp3826;
  assign tmp3826 = 1'b1;
  wire tmp3827;
  assign tmp3827 = ~pi5;
  wire tmp3828;
  assign tmp3828 = ~pi6;
  wire tmp3829;
  assign tmp3829 = (tmp3826 & tmp3827) | (tmp3826 & tmp3828) | (tmp3827 & tmp3828);
  wire tmp3830;
  assign tmp3830 = (tmp3821 & tmp3825) | (tmp3821 & tmp3829) | (tmp3825 & tmp3829);
  wire tmp3831;
  assign tmp3831 = 1'b1;
  wire tmp3832;
  assign tmp3832 = 1'b1;
  wire tmp3833;
  assign tmp3833 = 1'b1;
  wire tmp3834;
  assign tmp3834 = (tmp3831 & tmp3832) | (tmp3831 & tmp3833) | (tmp3832 & tmp3833);
  wire tmp3835;
  assign tmp3835 = 1'b1;
  wire tmp3836;
  assign tmp3836 = ~pi5;
  wire tmp3837;
  assign tmp3837 = ~pi6;
  wire tmp3838;
  assign tmp3838 = (tmp3835 & tmp3836) | (tmp3835 & tmp3837) | (tmp3836 & tmp3837);
  wire tmp3839;
  assign tmp3839 = 1'b1;
  wire tmp3840;
  assign tmp3840 = ~pi6;
  wire tmp3841;
  assign tmp3841 = ~pi7;
  wire tmp3842;
  assign tmp3842 = (tmp3839 & tmp3840) | (tmp3839 & tmp3841) | (tmp3840 & tmp3841);
  wire tmp3843;
  assign tmp3843 = (tmp3834 & tmp3838) | (tmp3834 & tmp3842) | (tmp3838 & tmp3842);
  wire tmp3844;
  assign tmp3844 = (tmp3817 & tmp3830) | (tmp3817 & tmp3843) | (tmp3830 & tmp3843);
  wire tmp3845;
  assign tmp3845 = 1'b0;
  wire tmp3846;
  assign tmp3846 = 1'b1;
  wire tmp3847;
  assign tmp3847 = 1'b0;
  wire tmp3848;
  assign tmp3848 = (tmp3845 & tmp3846) | (tmp3845 & tmp3847) | (tmp3846 & tmp3847);
  wire tmp3849;
  assign tmp3849 = 1'b1;
  wire tmp3850;
  assign tmp3850 = 1'b1;
  wire tmp3851;
  assign tmp3851 = 1'b1;
  wire tmp3852;
  assign tmp3852 = (tmp3849 & tmp3850) | (tmp3849 & tmp3851) | (tmp3850 & tmp3851);
  wire tmp3853;
  assign tmp3853 = 1'b0;
  wire tmp3854;
  assign tmp3854 = 1'b1;
  wire tmp3855;
  assign tmp3855 = 1'b0;
  wire tmp3856;
  assign tmp3856 = (tmp3853 & tmp3854) | (tmp3853 & tmp3855) | (tmp3854 & tmp3855);
  wire tmp3857;
  assign tmp3857 = (tmp3848 & tmp3852) | (tmp3848 & tmp3856) | (tmp3852 & tmp3856);
  wire tmp3858;
  assign tmp3858 = 1'b1;
  wire tmp3859;
  assign tmp3859 = 1'b1;
  wire tmp3860;
  assign tmp3860 = 1'b1;
  wire tmp3861;
  assign tmp3861 = (tmp3858 & tmp3859) | (tmp3858 & tmp3860) | (tmp3859 & tmp3860);
  wire tmp3862;
  assign tmp3862 = 1'b1;
  wire tmp3863;
  assign tmp3863 = ~pi5;
  wire tmp3864;
  assign tmp3864 = ~pi6;
  wire tmp3865;
  assign tmp3865 = (tmp3862 & tmp3863) | (tmp3862 & tmp3864) | (tmp3863 & tmp3864);
  wire tmp3866;
  assign tmp3866 = 1'b1;
  wire tmp3867;
  assign tmp3867 = ~pi6;
  wire tmp3868;
  assign tmp3868 = ~pi7;
  wire tmp3869;
  assign tmp3869 = (tmp3866 & tmp3867) | (tmp3866 & tmp3868) | (tmp3867 & tmp3868);
  wire tmp3870;
  assign tmp3870 = (tmp3861 & tmp3865) | (tmp3861 & tmp3869) | (tmp3865 & tmp3869);
  wire tmp3871;
  assign tmp3871 = 1'b0;
  wire tmp3872;
  assign tmp3872 = 1'b1;
  wire tmp3873;
  assign tmp3873 = 1'b0;
  wire tmp3874;
  assign tmp3874 = (tmp3871 & tmp3872) | (tmp3871 & tmp3873) | (tmp3872 & tmp3873);
  wire tmp3875;
  assign tmp3875 = 1'b1;
  wire tmp3876;
  assign tmp3876 = ~pi6;
  wire tmp3877;
  assign tmp3877 = ~pi7;
  wire tmp3878;
  assign tmp3878 = (tmp3875 & tmp3876) | (tmp3875 & tmp3877) | (tmp3876 & tmp3877);
  wire tmp3879;
  assign tmp3879 = 1'b0;
  wire tmp3880;
  assign tmp3880 = ~pi7;
  wire tmp3881;
  assign tmp3881 = 1'b0;
  wire tmp3882;
  assign tmp3882 = (tmp3879 & tmp3880) | (tmp3879 & tmp3881) | (tmp3880 & tmp3881);
  wire tmp3883;
  assign tmp3883 = (tmp3874 & tmp3878) | (tmp3874 & tmp3882) | (tmp3878 & tmp3882);
  wire tmp3884;
  assign tmp3884 = (tmp3857 & tmp3870) | (tmp3857 & tmp3883) | (tmp3870 & tmp3883);
  wire tmp3885;
  assign tmp3885 = (tmp3804 & tmp3844) | (tmp3804 & tmp3884) | (tmp3844 & tmp3884);
  wire tmp3886;
  assign tmp3886 = 1'b0;
  wire tmp3887;
  assign tmp3887 = 1'b0;
  wire tmp3888;
  assign tmp3888 = 1'b0;
  wire tmp3889;
  assign tmp3889 = (tmp3886 & tmp3887) | (tmp3886 & tmp3888) | (tmp3887 & tmp3888);
  wire tmp3890;
  assign tmp3890 = 1'b0;
  wire tmp3891;
  assign tmp3891 = 1'b1;
  wire tmp3892;
  assign tmp3892 = 1'b0;
  wire tmp3893;
  assign tmp3893 = (tmp3890 & tmp3891) | (tmp3890 & tmp3892) | (tmp3891 & tmp3892);
  wire tmp3894;
  assign tmp3894 = 1'b0;
  wire tmp3895;
  assign tmp3895 = 1'b0;
  wire tmp3896;
  assign tmp3896 = 1'b0;
  wire tmp3897;
  assign tmp3897 = (tmp3894 & tmp3895) | (tmp3894 & tmp3896) | (tmp3895 & tmp3896);
  wire tmp3898;
  assign tmp3898 = (tmp3889 & tmp3893) | (tmp3889 & tmp3897) | (tmp3893 & tmp3897);
  wire tmp3899;
  assign tmp3899 = 1'b0;
  wire tmp3900;
  assign tmp3900 = 1'b1;
  wire tmp3901;
  assign tmp3901 = 1'b0;
  wire tmp3902;
  assign tmp3902 = (tmp3899 & tmp3900) | (tmp3899 & tmp3901) | (tmp3900 & tmp3901);
  wire tmp3903;
  assign tmp3903 = 1'b1;
  wire tmp3904;
  assign tmp3904 = 1'b1;
  wire tmp3905;
  assign tmp3905 = 1'b1;
  wire tmp3906;
  assign tmp3906 = (tmp3903 & tmp3904) | (tmp3903 & tmp3905) | (tmp3904 & tmp3905);
  wire tmp3907;
  assign tmp3907 = 1'b0;
  wire tmp3908;
  assign tmp3908 = 1'b1;
  wire tmp3909;
  assign tmp3909 = 1'b0;
  wire tmp3910;
  assign tmp3910 = (tmp3907 & tmp3908) | (tmp3907 & tmp3909) | (tmp3908 & tmp3909);
  wire tmp3911;
  assign tmp3911 = (tmp3902 & tmp3906) | (tmp3902 & tmp3910) | (tmp3906 & tmp3910);
  wire tmp3912;
  assign tmp3912 = 1'b0;
  wire tmp3913;
  assign tmp3913 = 1'b0;
  wire tmp3914;
  assign tmp3914 = 1'b0;
  wire tmp3915;
  assign tmp3915 = (tmp3912 & tmp3913) | (tmp3912 & tmp3914) | (tmp3913 & tmp3914);
  wire tmp3916;
  assign tmp3916 = 1'b0;
  wire tmp3917;
  assign tmp3917 = 1'b1;
  wire tmp3918;
  assign tmp3918 = 1'b0;
  wire tmp3919;
  assign tmp3919 = (tmp3916 & tmp3917) | (tmp3916 & tmp3918) | (tmp3917 & tmp3918);
  wire tmp3920;
  assign tmp3920 = 1'b0;
  wire tmp3921;
  assign tmp3921 = 1'b0;
  wire tmp3922;
  assign tmp3922 = 1'b0;
  wire tmp3923;
  assign tmp3923 = (tmp3920 & tmp3921) | (tmp3920 & tmp3922) | (tmp3921 & tmp3922);
  wire tmp3924;
  assign tmp3924 = (tmp3915 & tmp3919) | (tmp3915 & tmp3923) | (tmp3919 & tmp3923);
  wire tmp3925;
  assign tmp3925 = (tmp3898 & tmp3911) | (tmp3898 & tmp3924) | (tmp3911 & tmp3924);
  wire tmp3926;
  assign tmp3926 = 1'b0;
  wire tmp3927;
  assign tmp3927 = 1'b1;
  wire tmp3928;
  assign tmp3928 = 1'b0;
  wire tmp3929;
  assign tmp3929 = (tmp3926 & tmp3927) | (tmp3926 & tmp3928) | (tmp3927 & tmp3928);
  wire tmp3930;
  assign tmp3930 = 1'b1;
  wire tmp3931;
  assign tmp3931 = 1'b1;
  wire tmp3932;
  assign tmp3932 = 1'b1;
  wire tmp3933;
  assign tmp3933 = (tmp3930 & tmp3931) | (tmp3930 & tmp3932) | (tmp3931 & tmp3932);
  wire tmp3934;
  assign tmp3934 = 1'b0;
  wire tmp3935;
  assign tmp3935 = 1'b1;
  wire tmp3936;
  assign tmp3936 = 1'b0;
  wire tmp3937;
  assign tmp3937 = (tmp3934 & tmp3935) | (tmp3934 & tmp3936) | (tmp3935 & tmp3936);
  wire tmp3938;
  assign tmp3938 = (tmp3929 & tmp3933) | (tmp3929 & tmp3937) | (tmp3933 & tmp3937);
  wire tmp3939;
  assign tmp3939 = 1'b1;
  wire tmp3940;
  assign tmp3940 = 1'b1;
  wire tmp3941;
  assign tmp3941 = 1'b1;
  wire tmp3942;
  assign tmp3942 = (tmp3939 & tmp3940) | (tmp3939 & tmp3941) | (tmp3940 & tmp3941);
  wire tmp3943;
  assign tmp3943 = 1'b1;
  wire tmp3944;
  assign tmp3944 = ~pi5;
  wire tmp3945;
  assign tmp3945 = ~pi6;
  wire tmp3946;
  assign tmp3946 = (tmp3943 & tmp3944) | (tmp3943 & tmp3945) | (tmp3944 & tmp3945);
  wire tmp3947;
  assign tmp3947 = 1'b1;
  wire tmp3948;
  assign tmp3948 = ~pi6;
  wire tmp3949;
  assign tmp3949 = ~pi7;
  wire tmp3950;
  assign tmp3950 = (tmp3947 & tmp3948) | (tmp3947 & tmp3949) | (tmp3948 & tmp3949);
  wire tmp3951;
  assign tmp3951 = (tmp3942 & tmp3946) | (tmp3942 & tmp3950) | (tmp3946 & tmp3950);
  wire tmp3952;
  assign tmp3952 = 1'b0;
  wire tmp3953;
  assign tmp3953 = 1'b1;
  wire tmp3954;
  assign tmp3954 = 1'b0;
  wire tmp3955;
  assign tmp3955 = (tmp3952 & tmp3953) | (tmp3952 & tmp3954) | (tmp3953 & tmp3954);
  wire tmp3956;
  assign tmp3956 = 1'b1;
  wire tmp3957;
  assign tmp3957 = ~pi6;
  wire tmp3958;
  assign tmp3958 = ~pi7;
  wire tmp3959;
  assign tmp3959 = (tmp3956 & tmp3957) | (tmp3956 & tmp3958) | (tmp3957 & tmp3958);
  wire tmp3960;
  assign tmp3960 = 1'b0;
  wire tmp3961;
  assign tmp3961 = ~pi7;
  wire tmp3962;
  assign tmp3962 = 1'b0;
  wire tmp3963;
  assign tmp3963 = (tmp3960 & tmp3961) | (tmp3960 & tmp3962) | (tmp3961 & tmp3962);
  wire tmp3964;
  assign tmp3964 = (tmp3955 & tmp3959) | (tmp3955 & tmp3963) | (tmp3959 & tmp3963);
  wire tmp3965;
  assign tmp3965 = (tmp3938 & tmp3951) | (tmp3938 & tmp3964) | (tmp3951 & tmp3964);
  wire tmp3966;
  assign tmp3966 = 1'b0;
  wire tmp3967;
  assign tmp3967 = 1'b0;
  wire tmp3968;
  assign tmp3968 = 1'b0;
  wire tmp3969;
  assign tmp3969 = (tmp3966 & tmp3967) | (tmp3966 & tmp3968) | (tmp3967 & tmp3968);
  wire tmp3970;
  assign tmp3970 = 1'b0;
  wire tmp3971;
  assign tmp3971 = 1'b1;
  wire tmp3972;
  assign tmp3972 = 1'b0;
  wire tmp3973;
  assign tmp3973 = (tmp3970 & tmp3971) | (tmp3970 & tmp3972) | (tmp3971 & tmp3972);
  wire tmp3974;
  assign tmp3974 = 1'b0;
  wire tmp3975;
  assign tmp3975 = 1'b0;
  wire tmp3976;
  assign tmp3976 = 1'b0;
  wire tmp3977;
  assign tmp3977 = (tmp3974 & tmp3975) | (tmp3974 & tmp3976) | (tmp3975 & tmp3976);
  wire tmp3978;
  assign tmp3978 = (tmp3969 & tmp3973) | (tmp3969 & tmp3977) | (tmp3973 & tmp3977);
  wire tmp3979;
  assign tmp3979 = 1'b0;
  wire tmp3980;
  assign tmp3980 = 1'b1;
  wire tmp3981;
  assign tmp3981 = 1'b0;
  wire tmp3982;
  assign tmp3982 = (tmp3979 & tmp3980) | (tmp3979 & tmp3981) | (tmp3980 & tmp3981);
  wire tmp3983;
  assign tmp3983 = 1'b1;
  wire tmp3984;
  assign tmp3984 = ~pi6;
  wire tmp3985;
  assign tmp3985 = ~pi7;
  wire tmp3986;
  assign tmp3986 = (tmp3983 & tmp3984) | (tmp3983 & tmp3985) | (tmp3984 & tmp3985);
  wire tmp3987;
  assign tmp3987 = 1'b0;
  wire tmp3988;
  assign tmp3988 = ~pi7;
  wire tmp3989;
  assign tmp3989 = 1'b0;
  wire tmp3990;
  assign tmp3990 = (tmp3987 & tmp3988) | (tmp3987 & tmp3989) | (tmp3988 & tmp3989);
  wire tmp3991;
  assign tmp3991 = (tmp3982 & tmp3986) | (tmp3982 & tmp3990) | (tmp3986 & tmp3990);
  wire tmp3992;
  assign tmp3992 = 1'b0;
  wire tmp3993;
  assign tmp3993 = 1'b0;
  wire tmp3994;
  assign tmp3994 = 1'b0;
  wire tmp3995;
  assign tmp3995 = (tmp3992 & tmp3993) | (tmp3992 & tmp3994) | (tmp3993 & tmp3994);
  wire tmp3996;
  assign tmp3996 = 1'b0;
  wire tmp3997;
  assign tmp3997 = ~pi7;
  wire tmp3998;
  assign tmp3998 = 1'b0;
  wire tmp3999;
  assign tmp3999 = (tmp3996 & tmp3997) | (tmp3996 & tmp3998) | (tmp3997 & tmp3998);
  wire tmp4000;
  assign tmp4000 = 1'b0;
  wire tmp4001;
  assign tmp4001 = 1'b0;
  wire tmp4002;
  assign tmp4002 = 1'b0;
  wire tmp4003;
  assign tmp4003 = (tmp4000 & tmp4001) | (tmp4000 & tmp4002) | (tmp4001 & tmp4002);
  wire tmp4004;
  assign tmp4004 = (tmp3995 & tmp3999) | (tmp3995 & tmp4003) | (tmp3999 & tmp4003);
  wire tmp4005;
  assign tmp4005 = (tmp3978 & tmp3991) | (tmp3978 & tmp4004) | (tmp3991 & tmp4004);
  wire tmp4006;
  assign tmp4006 = (tmp3925 & tmp3965) | (tmp3925 & tmp4005) | (tmp3965 & tmp4005);
  wire tmp4007;
  assign tmp4007 = (tmp3764 & tmp3885) | (tmp3764 & tmp4006) | (tmp3885 & tmp4006);
  wire tmp4008;
  assign tmp4008 = 1'b0;
  wire tmp4009;
  assign tmp4009 = 1'b0;
  wire tmp4010;
  assign tmp4010 = 1'b0;
  wire tmp4011;
  assign tmp4011 = (tmp4008 & tmp4009) | (tmp4008 & tmp4010) | (tmp4009 & tmp4010);
  wire tmp4012;
  assign tmp4012 = 1'b0;
  wire tmp4013;
  assign tmp4013 = 1'b0;
  wire tmp4014;
  assign tmp4014 = 1'b0;
  wire tmp4015;
  assign tmp4015 = (tmp4012 & tmp4013) | (tmp4012 & tmp4014) | (tmp4013 & tmp4014);
  wire tmp4016;
  assign tmp4016 = 1'b0;
  wire tmp4017;
  assign tmp4017 = 1'b0;
  wire tmp4018;
  assign tmp4018 = 1'b0;
  wire tmp4019;
  assign tmp4019 = (tmp4016 & tmp4017) | (tmp4016 & tmp4018) | (tmp4017 & tmp4018);
  wire tmp4020;
  assign tmp4020 = (tmp4011 & tmp4015) | (tmp4011 & tmp4019) | (tmp4015 & tmp4019);
  wire tmp4021;
  assign tmp4021 = 1'b0;
  wire tmp4022;
  assign tmp4022 = 1'b0;
  wire tmp4023;
  assign tmp4023 = 1'b0;
  wire tmp4024;
  assign tmp4024 = (tmp4021 & tmp4022) | (tmp4021 & tmp4023) | (tmp4022 & tmp4023);
  wire tmp4025;
  assign tmp4025 = 1'b0;
  wire tmp4026;
  assign tmp4026 = 1'b1;
  wire tmp4027;
  assign tmp4027 = 1'b0;
  wire tmp4028;
  assign tmp4028 = (tmp4025 & tmp4026) | (tmp4025 & tmp4027) | (tmp4026 & tmp4027);
  wire tmp4029;
  assign tmp4029 = 1'b0;
  wire tmp4030;
  assign tmp4030 = 1'b0;
  wire tmp4031;
  assign tmp4031 = 1'b0;
  wire tmp4032;
  assign tmp4032 = (tmp4029 & tmp4030) | (tmp4029 & tmp4031) | (tmp4030 & tmp4031);
  wire tmp4033;
  assign tmp4033 = (tmp4024 & tmp4028) | (tmp4024 & tmp4032) | (tmp4028 & tmp4032);
  wire tmp4034;
  assign tmp4034 = 1'b0;
  wire tmp4035;
  assign tmp4035 = 1'b0;
  wire tmp4036;
  assign tmp4036 = 1'b0;
  wire tmp4037;
  assign tmp4037 = (tmp4034 & tmp4035) | (tmp4034 & tmp4036) | (tmp4035 & tmp4036);
  wire tmp4038;
  assign tmp4038 = 1'b0;
  wire tmp4039;
  assign tmp4039 = 1'b0;
  wire tmp4040;
  assign tmp4040 = 1'b0;
  wire tmp4041;
  assign tmp4041 = (tmp4038 & tmp4039) | (tmp4038 & tmp4040) | (tmp4039 & tmp4040);
  wire tmp4042;
  assign tmp4042 = 1'b0;
  wire tmp4043;
  assign tmp4043 = 1'b0;
  wire tmp4044;
  assign tmp4044 = 1'b0;
  wire tmp4045;
  assign tmp4045 = (tmp4042 & tmp4043) | (tmp4042 & tmp4044) | (tmp4043 & tmp4044);
  wire tmp4046;
  assign tmp4046 = (tmp4037 & tmp4041) | (tmp4037 & tmp4045) | (tmp4041 & tmp4045);
  wire tmp4047;
  assign tmp4047 = (tmp4020 & tmp4033) | (tmp4020 & tmp4046) | (tmp4033 & tmp4046);
  wire tmp4048;
  assign tmp4048 = 1'b0;
  wire tmp4049;
  assign tmp4049 = 1'b0;
  wire tmp4050;
  assign tmp4050 = 1'b0;
  wire tmp4051;
  assign tmp4051 = (tmp4048 & tmp4049) | (tmp4048 & tmp4050) | (tmp4049 & tmp4050);
  wire tmp4052;
  assign tmp4052 = 1'b0;
  wire tmp4053;
  assign tmp4053 = 1'b1;
  wire tmp4054;
  assign tmp4054 = 1'b0;
  wire tmp4055;
  assign tmp4055 = (tmp4052 & tmp4053) | (tmp4052 & tmp4054) | (tmp4053 & tmp4054);
  wire tmp4056;
  assign tmp4056 = 1'b0;
  wire tmp4057;
  assign tmp4057 = 1'b0;
  wire tmp4058;
  assign tmp4058 = 1'b0;
  wire tmp4059;
  assign tmp4059 = (tmp4056 & tmp4057) | (tmp4056 & tmp4058) | (tmp4057 & tmp4058);
  wire tmp4060;
  assign tmp4060 = (tmp4051 & tmp4055) | (tmp4051 & tmp4059) | (tmp4055 & tmp4059);
  wire tmp4061;
  assign tmp4061 = 1'b0;
  wire tmp4062;
  assign tmp4062 = 1'b1;
  wire tmp4063;
  assign tmp4063 = 1'b0;
  wire tmp4064;
  assign tmp4064 = (tmp4061 & tmp4062) | (tmp4061 & tmp4063) | (tmp4062 & tmp4063);
  wire tmp4065;
  assign tmp4065 = 1'b1;
  wire tmp4066;
  assign tmp4066 = 1'b1;
  wire tmp4067;
  assign tmp4067 = 1'b1;
  wire tmp4068;
  assign tmp4068 = (tmp4065 & tmp4066) | (tmp4065 & tmp4067) | (tmp4066 & tmp4067);
  wire tmp4069;
  assign tmp4069 = 1'b0;
  wire tmp4070;
  assign tmp4070 = 1'b1;
  wire tmp4071;
  assign tmp4071 = 1'b0;
  wire tmp4072;
  assign tmp4072 = (tmp4069 & tmp4070) | (tmp4069 & tmp4071) | (tmp4070 & tmp4071);
  wire tmp4073;
  assign tmp4073 = (tmp4064 & tmp4068) | (tmp4064 & tmp4072) | (tmp4068 & tmp4072);
  wire tmp4074;
  assign tmp4074 = 1'b0;
  wire tmp4075;
  assign tmp4075 = 1'b0;
  wire tmp4076;
  assign tmp4076 = 1'b0;
  wire tmp4077;
  assign tmp4077 = (tmp4074 & tmp4075) | (tmp4074 & tmp4076) | (tmp4075 & tmp4076);
  wire tmp4078;
  assign tmp4078 = 1'b0;
  wire tmp4079;
  assign tmp4079 = 1'b1;
  wire tmp4080;
  assign tmp4080 = 1'b0;
  wire tmp4081;
  assign tmp4081 = (tmp4078 & tmp4079) | (tmp4078 & tmp4080) | (tmp4079 & tmp4080);
  wire tmp4082;
  assign tmp4082 = 1'b0;
  wire tmp4083;
  assign tmp4083 = 1'b0;
  wire tmp4084;
  assign tmp4084 = 1'b0;
  wire tmp4085;
  assign tmp4085 = (tmp4082 & tmp4083) | (tmp4082 & tmp4084) | (tmp4083 & tmp4084);
  wire tmp4086;
  assign tmp4086 = (tmp4077 & tmp4081) | (tmp4077 & tmp4085) | (tmp4081 & tmp4085);
  wire tmp4087;
  assign tmp4087 = (tmp4060 & tmp4073) | (tmp4060 & tmp4086) | (tmp4073 & tmp4086);
  wire tmp4088;
  assign tmp4088 = 1'b0;
  wire tmp4089;
  assign tmp4089 = 1'b0;
  wire tmp4090;
  assign tmp4090 = 1'b0;
  wire tmp4091;
  assign tmp4091 = (tmp4088 & tmp4089) | (tmp4088 & tmp4090) | (tmp4089 & tmp4090);
  wire tmp4092;
  assign tmp4092 = 1'b0;
  wire tmp4093;
  assign tmp4093 = 1'b0;
  wire tmp4094;
  assign tmp4094 = 1'b0;
  wire tmp4095;
  assign tmp4095 = (tmp4092 & tmp4093) | (tmp4092 & tmp4094) | (tmp4093 & tmp4094);
  wire tmp4096;
  assign tmp4096 = 1'b0;
  wire tmp4097;
  assign tmp4097 = 1'b0;
  wire tmp4098;
  assign tmp4098 = 1'b0;
  wire tmp4099;
  assign tmp4099 = (tmp4096 & tmp4097) | (tmp4096 & tmp4098) | (tmp4097 & tmp4098);
  wire tmp4100;
  assign tmp4100 = (tmp4091 & tmp4095) | (tmp4091 & tmp4099) | (tmp4095 & tmp4099);
  wire tmp4101;
  assign tmp4101 = 1'b0;
  wire tmp4102;
  assign tmp4102 = 1'b0;
  wire tmp4103;
  assign tmp4103 = 1'b0;
  wire tmp4104;
  assign tmp4104 = (tmp4101 & tmp4102) | (tmp4101 & tmp4103) | (tmp4102 & tmp4103);
  wire tmp4105;
  assign tmp4105 = 1'b0;
  wire tmp4106;
  assign tmp4106 = 1'b1;
  wire tmp4107;
  assign tmp4107 = 1'b0;
  wire tmp4108;
  assign tmp4108 = (tmp4105 & tmp4106) | (tmp4105 & tmp4107) | (tmp4106 & tmp4107);
  wire tmp4109;
  assign tmp4109 = 1'b0;
  wire tmp4110;
  assign tmp4110 = 1'b0;
  wire tmp4111;
  assign tmp4111 = 1'b0;
  wire tmp4112;
  assign tmp4112 = (tmp4109 & tmp4110) | (tmp4109 & tmp4111) | (tmp4110 & tmp4111);
  wire tmp4113;
  assign tmp4113 = (tmp4104 & tmp4108) | (tmp4104 & tmp4112) | (tmp4108 & tmp4112);
  wire tmp4114;
  assign tmp4114 = 1'b0;
  wire tmp4115;
  assign tmp4115 = 1'b0;
  wire tmp4116;
  assign tmp4116 = 1'b0;
  wire tmp4117;
  assign tmp4117 = (tmp4114 & tmp4115) | (tmp4114 & tmp4116) | (tmp4115 & tmp4116);
  wire tmp4118;
  assign tmp4118 = 1'b0;
  wire tmp4119;
  assign tmp4119 = 1'b0;
  wire tmp4120;
  assign tmp4120 = 1'b0;
  wire tmp4121;
  assign tmp4121 = (tmp4118 & tmp4119) | (tmp4118 & tmp4120) | (tmp4119 & tmp4120);
  wire tmp4122;
  assign tmp4122 = 1'b0;
  wire tmp4123;
  assign tmp4123 = 1'b0;
  wire tmp4124;
  assign tmp4124 = 1'b0;
  wire tmp4125;
  assign tmp4125 = (tmp4122 & tmp4123) | (tmp4122 & tmp4124) | (tmp4123 & tmp4124);
  wire tmp4126;
  assign tmp4126 = (tmp4117 & tmp4121) | (tmp4117 & tmp4125) | (tmp4121 & tmp4125);
  wire tmp4127;
  assign tmp4127 = (tmp4100 & tmp4113) | (tmp4100 & tmp4126) | (tmp4113 & tmp4126);
  wire tmp4128;
  assign tmp4128 = (tmp4047 & tmp4087) | (tmp4047 & tmp4127) | (tmp4087 & tmp4127);
  wire tmp4129;
  assign tmp4129 = 1'b0;
  wire tmp4130;
  assign tmp4130 = 1'b0;
  wire tmp4131;
  assign tmp4131 = 1'b0;
  wire tmp4132;
  assign tmp4132 = (tmp4129 & tmp4130) | (tmp4129 & tmp4131) | (tmp4130 & tmp4131);
  wire tmp4133;
  assign tmp4133 = 1'b0;
  wire tmp4134;
  assign tmp4134 = 1'b1;
  wire tmp4135;
  assign tmp4135 = 1'b0;
  wire tmp4136;
  assign tmp4136 = (tmp4133 & tmp4134) | (tmp4133 & tmp4135) | (tmp4134 & tmp4135);
  wire tmp4137;
  assign tmp4137 = 1'b0;
  wire tmp4138;
  assign tmp4138 = 1'b0;
  wire tmp4139;
  assign tmp4139 = 1'b0;
  wire tmp4140;
  assign tmp4140 = (tmp4137 & tmp4138) | (tmp4137 & tmp4139) | (tmp4138 & tmp4139);
  wire tmp4141;
  assign tmp4141 = (tmp4132 & tmp4136) | (tmp4132 & tmp4140) | (tmp4136 & tmp4140);
  wire tmp4142;
  assign tmp4142 = 1'b0;
  wire tmp4143;
  assign tmp4143 = 1'b1;
  wire tmp4144;
  assign tmp4144 = 1'b0;
  wire tmp4145;
  assign tmp4145 = (tmp4142 & tmp4143) | (tmp4142 & tmp4144) | (tmp4143 & tmp4144);
  wire tmp4146;
  assign tmp4146 = 1'b1;
  wire tmp4147;
  assign tmp4147 = 1'b1;
  wire tmp4148;
  assign tmp4148 = 1'b1;
  wire tmp4149;
  assign tmp4149 = (tmp4146 & tmp4147) | (tmp4146 & tmp4148) | (tmp4147 & tmp4148);
  wire tmp4150;
  assign tmp4150 = 1'b0;
  wire tmp4151;
  assign tmp4151 = 1'b1;
  wire tmp4152;
  assign tmp4152 = 1'b0;
  wire tmp4153;
  assign tmp4153 = (tmp4150 & tmp4151) | (tmp4150 & tmp4152) | (tmp4151 & tmp4152);
  wire tmp4154;
  assign tmp4154 = (tmp4145 & tmp4149) | (tmp4145 & tmp4153) | (tmp4149 & tmp4153);
  wire tmp4155;
  assign tmp4155 = 1'b0;
  wire tmp4156;
  assign tmp4156 = 1'b0;
  wire tmp4157;
  assign tmp4157 = 1'b0;
  wire tmp4158;
  assign tmp4158 = (tmp4155 & tmp4156) | (tmp4155 & tmp4157) | (tmp4156 & tmp4157);
  wire tmp4159;
  assign tmp4159 = 1'b0;
  wire tmp4160;
  assign tmp4160 = 1'b1;
  wire tmp4161;
  assign tmp4161 = 1'b0;
  wire tmp4162;
  assign tmp4162 = (tmp4159 & tmp4160) | (tmp4159 & tmp4161) | (tmp4160 & tmp4161);
  wire tmp4163;
  assign tmp4163 = 1'b0;
  wire tmp4164;
  assign tmp4164 = 1'b0;
  wire tmp4165;
  assign tmp4165 = 1'b0;
  wire tmp4166;
  assign tmp4166 = (tmp4163 & tmp4164) | (tmp4163 & tmp4165) | (tmp4164 & tmp4165);
  wire tmp4167;
  assign tmp4167 = (tmp4158 & tmp4162) | (tmp4158 & tmp4166) | (tmp4162 & tmp4166);
  wire tmp4168;
  assign tmp4168 = (tmp4141 & tmp4154) | (tmp4141 & tmp4167) | (tmp4154 & tmp4167);
  wire tmp4169;
  assign tmp4169 = 1'b0;
  wire tmp4170;
  assign tmp4170 = 1'b1;
  wire tmp4171;
  assign tmp4171 = 1'b0;
  wire tmp4172;
  assign tmp4172 = (tmp4169 & tmp4170) | (tmp4169 & tmp4171) | (tmp4170 & tmp4171);
  wire tmp4173;
  assign tmp4173 = 1'b1;
  wire tmp4174;
  assign tmp4174 = 1'b1;
  wire tmp4175;
  assign tmp4175 = 1'b1;
  wire tmp4176;
  assign tmp4176 = (tmp4173 & tmp4174) | (tmp4173 & tmp4175) | (tmp4174 & tmp4175);
  wire tmp4177;
  assign tmp4177 = 1'b0;
  wire tmp4178;
  assign tmp4178 = 1'b1;
  wire tmp4179;
  assign tmp4179 = 1'b0;
  wire tmp4180;
  assign tmp4180 = (tmp4177 & tmp4178) | (tmp4177 & tmp4179) | (tmp4178 & tmp4179);
  wire tmp4181;
  assign tmp4181 = (tmp4172 & tmp4176) | (tmp4172 & tmp4180) | (tmp4176 & tmp4180);
  wire tmp4182;
  assign tmp4182 = 1'b1;
  wire tmp4183;
  assign tmp4183 = 1'b1;
  wire tmp4184;
  assign tmp4184 = 1'b1;
  wire tmp4185;
  assign tmp4185 = (tmp4182 & tmp4183) | (tmp4182 & tmp4184) | (tmp4183 & tmp4184);
  wire tmp4186;
  assign tmp4186 = 1'b1;
  wire tmp4187;
  assign tmp4187 = ~pi5;
  wire tmp4188;
  assign tmp4188 = ~pi6;
  wire tmp4189;
  assign tmp4189 = (tmp4186 & tmp4187) | (tmp4186 & tmp4188) | (tmp4187 & tmp4188);
  wire tmp4190;
  assign tmp4190 = 1'b1;
  wire tmp4191;
  assign tmp4191 = ~pi6;
  wire tmp4192;
  assign tmp4192 = ~pi7;
  wire tmp4193;
  assign tmp4193 = (tmp4190 & tmp4191) | (tmp4190 & tmp4192) | (tmp4191 & tmp4192);
  wire tmp4194;
  assign tmp4194 = (tmp4185 & tmp4189) | (tmp4185 & tmp4193) | (tmp4189 & tmp4193);
  wire tmp4195;
  assign tmp4195 = 1'b0;
  wire tmp4196;
  assign tmp4196 = 1'b1;
  wire tmp4197;
  assign tmp4197 = 1'b0;
  wire tmp4198;
  assign tmp4198 = (tmp4195 & tmp4196) | (tmp4195 & tmp4197) | (tmp4196 & tmp4197);
  wire tmp4199;
  assign tmp4199 = 1'b1;
  wire tmp4200;
  assign tmp4200 = ~pi6;
  wire tmp4201;
  assign tmp4201 = ~pi7;
  wire tmp4202;
  assign tmp4202 = (tmp4199 & tmp4200) | (tmp4199 & tmp4201) | (tmp4200 & tmp4201);
  wire tmp4203;
  assign tmp4203 = 1'b0;
  wire tmp4204;
  assign tmp4204 = ~pi7;
  wire tmp4205;
  assign tmp4205 = 1'b0;
  wire tmp4206;
  assign tmp4206 = (tmp4203 & tmp4204) | (tmp4203 & tmp4205) | (tmp4204 & tmp4205);
  wire tmp4207;
  assign tmp4207 = (tmp4198 & tmp4202) | (tmp4198 & tmp4206) | (tmp4202 & tmp4206);
  wire tmp4208;
  assign tmp4208 = (tmp4181 & tmp4194) | (tmp4181 & tmp4207) | (tmp4194 & tmp4207);
  wire tmp4209;
  assign tmp4209 = 1'b0;
  wire tmp4210;
  assign tmp4210 = 1'b0;
  wire tmp4211;
  assign tmp4211 = 1'b0;
  wire tmp4212;
  assign tmp4212 = (tmp4209 & tmp4210) | (tmp4209 & tmp4211) | (tmp4210 & tmp4211);
  wire tmp4213;
  assign tmp4213 = 1'b0;
  wire tmp4214;
  assign tmp4214 = 1'b1;
  wire tmp4215;
  assign tmp4215 = 1'b0;
  wire tmp4216;
  assign tmp4216 = (tmp4213 & tmp4214) | (tmp4213 & tmp4215) | (tmp4214 & tmp4215);
  wire tmp4217;
  assign tmp4217 = 1'b0;
  wire tmp4218;
  assign tmp4218 = 1'b0;
  wire tmp4219;
  assign tmp4219 = 1'b0;
  wire tmp4220;
  assign tmp4220 = (tmp4217 & tmp4218) | (tmp4217 & tmp4219) | (tmp4218 & tmp4219);
  wire tmp4221;
  assign tmp4221 = (tmp4212 & tmp4216) | (tmp4212 & tmp4220) | (tmp4216 & tmp4220);
  wire tmp4222;
  assign tmp4222 = 1'b0;
  wire tmp4223;
  assign tmp4223 = 1'b1;
  wire tmp4224;
  assign tmp4224 = 1'b0;
  wire tmp4225;
  assign tmp4225 = (tmp4222 & tmp4223) | (tmp4222 & tmp4224) | (tmp4223 & tmp4224);
  wire tmp4226;
  assign tmp4226 = 1'b1;
  wire tmp4227;
  assign tmp4227 = ~pi6;
  wire tmp4228;
  assign tmp4228 = ~pi7;
  wire tmp4229;
  assign tmp4229 = (tmp4226 & tmp4227) | (tmp4226 & tmp4228) | (tmp4227 & tmp4228);
  wire tmp4230;
  assign tmp4230 = 1'b0;
  wire tmp4231;
  assign tmp4231 = ~pi7;
  wire tmp4232;
  assign tmp4232 = 1'b0;
  wire tmp4233;
  assign tmp4233 = (tmp4230 & tmp4231) | (tmp4230 & tmp4232) | (tmp4231 & tmp4232);
  wire tmp4234;
  assign tmp4234 = (tmp4225 & tmp4229) | (tmp4225 & tmp4233) | (tmp4229 & tmp4233);
  wire tmp4235;
  assign tmp4235 = 1'b0;
  wire tmp4236;
  assign tmp4236 = 1'b0;
  wire tmp4237;
  assign tmp4237 = 1'b0;
  wire tmp4238;
  assign tmp4238 = (tmp4235 & tmp4236) | (tmp4235 & tmp4237) | (tmp4236 & tmp4237);
  wire tmp4239;
  assign tmp4239 = 1'b0;
  wire tmp4240;
  assign tmp4240 = ~pi7;
  wire tmp4241;
  assign tmp4241 = 1'b0;
  wire tmp4242;
  assign tmp4242 = (tmp4239 & tmp4240) | (tmp4239 & tmp4241) | (tmp4240 & tmp4241);
  wire tmp4243;
  assign tmp4243 = 1'b0;
  wire tmp4244;
  assign tmp4244 = 1'b0;
  wire tmp4245;
  assign tmp4245 = 1'b0;
  wire tmp4246;
  assign tmp4246 = (tmp4243 & tmp4244) | (tmp4243 & tmp4245) | (tmp4244 & tmp4245);
  wire tmp4247;
  assign tmp4247 = (tmp4238 & tmp4242) | (tmp4238 & tmp4246) | (tmp4242 & tmp4246);
  wire tmp4248;
  assign tmp4248 = (tmp4221 & tmp4234) | (tmp4221 & tmp4247) | (tmp4234 & tmp4247);
  wire tmp4249;
  assign tmp4249 = (tmp4168 & tmp4208) | (tmp4168 & tmp4248) | (tmp4208 & tmp4248);
  wire tmp4250;
  assign tmp4250 = 1'b0;
  wire tmp4251;
  assign tmp4251 = 1'b0;
  wire tmp4252;
  assign tmp4252 = 1'b0;
  wire tmp4253;
  assign tmp4253 = (tmp4250 & tmp4251) | (tmp4250 & tmp4252) | (tmp4251 & tmp4252);
  wire tmp4254;
  assign tmp4254 = 1'b0;
  wire tmp4255;
  assign tmp4255 = 1'b0;
  wire tmp4256;
  assign tmp4256 = 1'b0;
  wire tmp4257;
  assign tmp4257 = (tmp4254 & tmp4255) | (tmp4254 & tmp4256) | (tmp4255 & tmp4256);
  wire tmp4258;
  assign tmp4258 = 1'b0;
  wire tmp4259;
  assign tmp4259 = 1'b0;
  wire tmp4260;
  assign tmp4260 = 1'b0;
  wire tmp4261;
  assign tmp4261 = (tmp4258 & tmp4259) | (tmp4258 & tmp4260) | (tmp4259 & tmp4260);
  wire tmp4262;
  assign tmp4262 = (tmp4253 & tmp4257) | (tmp4253 & tmp4261) | (tmp4257 & tmp4261);
  wire tmp4263;
  assign tmp4263 = 1'b0;
  wire tmp4264;
  assign tmp4264 = 1'b0;
  wire tmp4265;
  assign tmp4265 = 1'b0;
  wire tmp4266;
  assign tmp4266 = (tmp4263 & tmp4264) | (tmp4263 & tmp4265) | (tmp4264 & tmp4265);
  wire tmp4267;
  assign tmp4267 = 1'b0;
  wire tmp4268;
  assign tmp4268 = 1'b1;
  wire tmp4269;
  assign tmp4269 = 1'b0;
  wire tmp4270;
  assign tmp4270 = (tmp4267 & tmp4268) | (tmp4267 & tmp4269) | (tmp4268 & tmp4269);
  wire tmp4271;
  assign tmp4271 = 1'b0;
  wire tmp4272;
  assign tmp4272 = 1'b0;
  wire tmp4273;
  assign tmp4273 = 1'b0;
  wire tmp4274;
  assign tmp4274 = (tmp4271 & tmp4272) | (tmp4271 & tmp4273) | (tmp4272 & tmp4273);
  wire tmp4275;
  assign tmp4275 = (tmp4266 & tmp4270) | (tmp4266 & tmp4274) | (tmp4270 & tmp4274);
  wire tmp4276;
  assign tmp4276 = 1'b0;
  wire tmp4277;
  assign tmp4277 = 1'b0;
  wire tmp4278;
  assign tmp4278 = 1'b0;
  wire tmp4279;
  assign tmp4279 = (tmp4276 & tmp4277) | (tmp4276 & tmp4278) | (tmp4277 & tmp4278);
  wire tmp4280;
  assign tmp4280 = 1'b0;
  wire tmp4281;
  assign tmp4281 = 1'b0;
  wire tmp4282;
  assign tmp4282 = 1'b0;
  wire tmp4283;
  assign tmp4283 = (tmp4280 & tmp4281) | (tmp4280 & tmp4282) | (tmp4281 & tmp4282);
  wire tmp4284;
  assign tmp4284 = 1'b0;
  wire tmp4285;
  assign tmp4285 = 1'b0;
  wire tmp4286;
  assign tmp4286 = 1'b0;
  wire tmp4287;
  assign tmp4287 = (tmp4284 & tmp4285) | (tmp4284 & tmp4286) | (tmp4285 & tmp4286);
  wire tmp4288;
  assign tmp4288 = (tmp4279 & tmp4283) | (tmp4279 & tmp4287) | (tmp4283 & tmp4287);
  wire tmp4289;
  assign tmp4289 = (tmp4262 & tmp4275) | (tmp4262 & tmp4288) | (tmp4275 & tmp4288);
  wire tmp4290;
  assign tmp4290 = 1'b0;
  wire tmp4291;
  assign tmp4291 = 1'b0;
  wire tmp4292;
  assign tmp4292 = 1'b0;
  wire tmp4293;
  assign tmp4293 = (tmp4290 & tmp4291) | (tmp4290 & tmp4292) | (tmp4291 & tmp4292);
  wire tmp4294;
  assign tmp4294 = 1'b0;
  wire tmp4295;
  assign tmp4295 = 1'b1;
  wire tmp4296;
  assign tmp4296 = 1'b0;
  wire tmp4297;
  assign tmp4297 = (tmp4294 & tmp4295) | (tmp4294 & tmp4296) | (tmp4295 & tmp4296);
  wire tmp4298;
  assign tmp4298 = 1'b0;
  wire tmp4299;
  assign tmp4299 = 1'b0;
  wire tmp4300;
  assign tmp4300 = 1'b0;
  wire tmp4301;
  assign tmp4301 = (tmp4298 & tmp4299) | (tmp4298 & tmp4300) | (tmp4299 & tmp4300);
  wire tmp4302;
  assign tmp4302 = (tmp4293 & tmp4297) | (tmp4293 & tmp4301) | (tmp4297 & tmp4301);
  wire tmp4303;
  assign tmp4303 = 1'b0;
  wire tmp4304;
  assign tmp4304 = 1'b1;
  wire tmp4305;
  assign tmp4305 = 1'b0;
  wire tmp4306;
  assign tmp4306 = (tmp4303 & tmp4304) | (tmp4303 & tmp4305) | (tmp4304 & tmp4305);
  wire tmp4307;
  assign tmp4307 = 1'b1;
  wire tmp4308;
  assign tmp4308 = ~pi6;
  wire tmp4309;
  assign tmp4309 = ~pi7;
  wire tmp4310;
  assign tmp4310 = (tmp4307 & tmp4308) | (tmp4307 & tmp4309) | (tmp4308 & tmp4309);
  wire tmp4311;
  assign tmp4311 = 1'b0;
  wire tmp4312;
  assign tmp4312 = ~pi7;
  wire tmp4313;
  assign tmp4313 = 1'b0;
  wire tmp4314;
  assign tmp4314 = (tmp4311 & tmp4312) | (tmp4311 & tmp4313) | (tmp4312 & tmp4313);
  wire tmp4315;
  assign tmp4315 = (tmp4306 & tmp4310) | (tmp4306 & tmp4314) | (tmp4310 & tmp4314);
  wire tmp4316;
  assign tmp4316 = 1'b0;
  wire tmp4317;
  assign tmp4317 = 1'b0;
  wire tmp4318;
  assign tmp4318 = 1'b0;
  wire tmp4319;
  assign tmp4319 = (tmp4316 & tmp4317) | (tmp4316 & tmp4318) | (tmp4317 & tmp4318);
  wire tmp4320;
  assign tmp4320 = 1'b0;
  wire tmp4321;
  assign tmp4321 = ~pi7;
  wire tmp4322;
  assign tmp4322 = 1'b0;
  wire tmp4323;
  assign tmp4323 = (tmp4320 & tmp4321) | (tmp4320 & tmp4322) | (tmp4321 & tmp4322);
  wire tmp4324;
  assign tmp4324 = 1'b0;
  wire tmp4325;
  assign tmp4325 = 1'b0;
  wire tmp4326;
  assign tmp4326 = 1'b0;
  wire tmp4327;
  assign tmp4327 = (tmp4324 & tmp4325) | (tmp4324 & tmp4326) | (tmp4325 & tmp4326);
  wire tmp4328;
  assign tmp4328 = (tmp4319 & tmp4323) | (tmp4319 & tmp4327) | (tmp4323 & tmp4327);
  wire tmp4329;
  assign tmp4329 = (tmp4302 & tmp4315) | (tmp4302 & tmp4328) | (tmp4315 & tmp4328);
  wire tmp4330;
  assign tmp4330 = 1'b0;
  wire tmp4331;
  assign tmp4331 = 1'b0;
  wire tmp4332;
  assign tmp4332 = 1'b0;
  wire tmp4333;
  assign tmp4333 = (tmp4330 & tmp4331) | (tmp4330 & tmp4332) | (tmp4331 & tmp4332);
  wire tmp4334;
  assign tmp4334 = 1'b0;
  wire tmp4335;
  assign tmp4335 = 1'b0;
  wire tmp4336;
  assign tmp4336 = 1'b0;
  wire tmp4337;
  assign tmp4337 = (tmp4334 & tmp4335) | (tmp4334 & tmp4336) | (tmp4335 & tmp4336);
  wire tmp4338;
  assign tmp4338 = 1'b0;
  wire tmp4339;
  assign tmp4339 = 1'b0;
  wire tmp4340;
  assign tmp4340 = 1'b0;
  wire tmp4341;
  assign tmp4341 = (tmp4338 & tmp4339) | (tmp4338 & tmp4340) | (tmp4339 & tmp4340);
  wire tmp4342;
  assign tmp4342 = (tmp4333 & tmp4337) | (tmp4333 & tmp4341) | (tmp4337 & tmp4341);
  wire tmp4343;
  assign tmp4343 = 1'b0;
  wire tmp4344;
  assign tmp4344 = 1'b0;
  wire tmp4345;
  assign tmp4345 = 1'b0;
  wire tmp4346;
  assign tmp4346 = (tmp4343 & tmp4344) | (tmp4343 & tmp4345) | (tmp4344 & tmp4345);
  wire tmp4347;
  assign tmp4347 = 1'b0;
  wire tmp4348;
  assign tmp4348 = ~pi7;
  wire tmp4349;
  assign tmp4349 = 1'b0;
  wire tmp4350;
  assign tmp4350 = (tmp4347 & tmp4348) | (tmp4347 & tmp4349) | (tmp4348 & tmp4349);
  wire tmp4351;
  assign tmp4351 = 1'b0;
  wire tmp4352;
  assign tmp4352 = 1'b0;
  wire tmp4353;
  assign tmp4353 = 1'b0;
  wire tmp4354;
  assign tmp4354 = (tmp4351 & tmp4352) | (tmp4351 & tmp4353) | (tmp4352 & tmp4353);
  wire tmp4355;
  assign tmp4355 = (tmp4346 & tmp4350) | (tmp4346 & tmp4354) | (tmp4350 & tmp4354);
  wire tmp4356;
  assign tmp4356 = 1'b0;
  wire tmp4357;
  assign tmp4357 = 1'b0;
  wire tmp4358;
  assign tmp4358 = 1'b0;
  wire tmp4359;
  assign tmp4359 = (tmp4356 & tmp4357) | (tmp4356 & tmp4358) | (tmp4357 & tmp4358);
  wire tmp4360;
  assign tmp4360 = 1'b0;
  wire tmp4361;
  assign tmp4361 = 1'b0;
  wire tmp4362;
  assign tmp4362 = 1'b0;
  wire tmp4363;
  assign tmp4363 = (tmp4360 & tmp4361) | (tmp4360 & tmp4362) | (tmp4361 & tmp4362);
  wire tmp4364;
  assign tmp4364 = 1'b0;
  wire tmp4365;
  assign tmp4365 = 1'b0;
  wire tmp4366;
  assign tmp4366 = 1'b0;
  wire tmp4367;
  assign tmp4367 = (tmp4364 & tmp4365) | (tmp4364 & tmp4366) | (tmp4365 & tmp4366);
  wire tmp4368;
  assign tmp4368 = (tmp4359 & tmp4363) | (tmp4359 & tmp4367) | (tmp4363 & tmp4367);
  wire tmp4369;
  assign tmp4369 = (tmp4342 & tmp4355) | (tmp4342 & tmp4368) | (tmp4355 & tmp4368);
  wire tmp4370;
  assign tmp4370 = (tmp4289 & tmp4329) | (tmp4289 & tmp4369) | (tmp4329 & tmp4369);
  wire tmp4371;
  assign tmp4371 = (tmp4128 & tmp4249) | (tmp4128 & tmp4370) | (tmp4249 & tmp4370);
  wire tmp4372;
  assign tmp4372 = (tmp3643 & tmp4007) | (tmp3643 & tmp4371) | (tmp4007 & tmp4371);
  wire tmp4373;
  assign tmp4373 = pi2;
  wire tmp4374;
  assign tmp4374 = pi3;
  wire tmp4375;
  assign tmp4375 = 1'b0;
  wire tmp4376;
  assign tmp4376 = (tmp4373 & tmp4374) | (tmp4373 & tmp4375) | (tmp4374 & tmp4375);
  wire tmp4377;
  assign tmp4377 = pi3;
  wire tmp4378;
  assign tmp4378 = 1'b1;
  wire tmp4379;
  assign tmp4379 = 1'b0;
  wire tmp4380;
  assign tmp4380 = (tmp4377 & tmp4378) | (tmp4377 & tmp4379) | (tmp4378 & tmp4379);
  wire tmp4381;
  assign tmp4381 = 1'b0;
  wire tmp4382;
  assign tmp4382 = 1'b0;
  wire tmp4383;
  assign tmp4383 = 1'b0;
  wire tmp4384;
  assign tmp4384 = (tmp4381 & tmp4382) | (tmp4381 & tmp4383) | (tmp4382 & tmp4383);
  wire tmp4385;
  assign tmp4385 = (tmp4376 & tmp4380) | (tmp4376 & tmp4384) | (tmp4380 & tmp4384);
  wire tmp4386;
  assign tmp4386 = pi3;
  wire tmp4387;
  assign tmp4387 = 1'b1;
  wire tmp4388;
  assign tmp4388 = 1'b0;
  wire tmp4389;
  assign tmp4389 = (tmp4386 & tmp4387) | (tmp4386 & tmp4388) | (tmp4387 & tmp4388);
  wire tmp4390;
  assign tmp4390 = 1'b1;
  wire tmp4391;
  assign tmp4391 = 1'b1;
  wire tmp4392;
  assign tmp4392 = 1'b1;
  wire tmp4393;
  assign tmp4393 = (tmp4390 & tmp4391) | (tmp4390 & tmp4392) | (tmp4391 & tmp4392);
  wire tmp4394;
  assign tmp4394 = 1'b0;
  wire tmp4395;
  assign tmp4395 = 1'b1;
  wire tmp4396;
  assign tmp4396 = 1'b0;
  wire tmp4397;
  assign tmp4397 = (tmp4394 & tmp4395) | (tmp4394 & tmp4396) | (tmp4395 & tmp4396);
  wire tmp4398;
  assign tmp4398 = (tmp4389 & tmp4393) | (tmp4389 & tmp4397) | (tmp4393 & tmp4397);
  wire tmp4399;
  assign tmp4399 = 1'b0;
  wire tmp4400;
  assign tmp4400 = 1'b0;
  wire tmp4401;
  assign tmp4401 = 1'b0;
  wire tmp4402;
  assign tmp4402 = (tmp4399 & tmp4400) | (tmp4399 & tmp4401) | (tmp4400 & tmp4401);
  wire tmp4403;
  assign tmp4403 = 1'b0;
  wire tmp4404;
  assign tmp4404 = 1'b1;
  wire tmp4405;
  assign tmp4405 = 1'b0;
  wire tmp4406;
  assign tmp4406 = (tmp4403 & tmp4404) | (tmp4403 & tmp4405) | (tmp4404 & tmp4405);
  wire tmp4407;
  assign tmp4407 = 1'b0;
  wire tmp4408;
  assign tmp4408 = 1'b0;
  wire tmp4409;
  assign tmp4409 = 1'b0;
  wire tmp4410;
  assign tmp4410 = (tmp4407 & tmp4408) | (tmp4407 & tmp4409) | (tmp4408 & tmp4409);
  wire tmp4411;
  assign tmp4411 = (tmp4402 & tmp4406) | (tmp4402 & tmp4410) | (tmp4406 & tmp4410);
  wire tmp4412;
  assign tmp4412 = (tmp4385 & tmp4398) | (tmp4385 & tmp4411) | (tmp4398 & tmp4411);
  wire tmp4413;
  assign tmp4413 = pi3;
  wire tmp4414;
  assign tmp4414 = 1'b1;
  wire tmp4415;
  assign tmp4415 = 1'b0;
  wire tmp4416;
  assign tmp4416 = (tmp4413 & tmp4414) | (tmp4413 & tmp4415) | (tmp4414 & tmp4415);
  wire tmp4417;
  assign tmp4417 = 1'b1;
  wire tmp4418;
  assign tmp4418 = 1'b1;
  wire tmp4419;
  assign tmp4419 = 1'b1;
  wire tmp4420;
  assign tmp4420 = (tmp4417 & tmp4418) | (tmp4417 & tmp4419) | (tmp4418 & tmp4419);
  wire tmp4421;
  assign tmp4421 = 1'b0;
  wire tmp4422;
  assign tmp4422 = 1'b1;
  wire tmp4423;
  assign tmp4423 = 1'b0;
  wire tmp4424;
  assign tmp4424 = (tmp4421 & tmp4422) | (tmp4421 & tmp4423) | (tmp4422 & tmp4423);
  wire tmp4425;
  assign tmp4425 = (tmp4416 & tmp4420) | (tmp4416 & tmp4424) | (tmp4420 & tmp4424);
  wire tmp4426;
  assign tmp4426 = 1'b1;
  wire tmp4427;
  assign tmp4427 = 1'b1;
  wire tmp4428;
  assign tmp4428 = 1'b1;
  wire tmp4429;
  assign tmp4429 = (tmp4426 & tmp4427) | (tmp4426 & tmp4428) | (tmp4427 & tmp4428);
  wire tmp4430;
  assign tmp4430 = 1'b1;
  wire tmp4431;
  assign tmp4431 = 1'b1;
  wire tmp4432;
  assign tmp4432 = 1'b1;
  wire tmp4433;
  assign tmp4433 = (tmp4430 & tmp4431) | (tmp4430 & tmp4432) | (tmp4431 & tmp4432);
  wire tmp4434;
  assign tmp4434 = 1'b1;
  wire tmp4435;
  assign tmp4435 = 1'b1;
  wire tmp4436;
  assign tmp4436 = 1'b1;
  wire tmp4437;
  assign tmp4437 = (tmp4434 & tmp4435) | (tmp4434 & tmp4436) | (tmp4435 & tmp4436);
  wire tmp4438;
  assign tmp4438 = (tmp4429 & tmp4433) | (tmp4429 & tmp4437) | (tmp4433 & tmp4437);
  wire tmp4439;
  assign tmp4439 = 1'b0;
  wire tmp4440;
  assign tmp4440 = 1'b1;
  wire tmp4441;
  assign tmp4441 = 1'b0;
  wire tmp4442;
  assign tmp4442 = (tmp4439 & tmp4440) | (tmp4439 & tmp4441) | (tmp4440 & tmp4441);
  wire tmp4443;
  assign tmp4443 = 1'b1;
  wire tmp4444;
  assign tmp4444 = 1'b1;
  wire tmp4445;
  assign tmp4445 = 1'b1;
  wire tmp4446;
  assign tmp4446 = (tmp4443 & tmp4444) | (tmp4443 & tmp4445) | (tmp4444 & tmp4445);
  wire tmp4447;
  assign tmp4447 = 1'b0;
  wire tmp4448;
  assign tmp4448 = 1'b1;
  wire tmp4449;
  assign tmp4449 = 1'b0;
  wire tmp4450;
  assign tmp4450 = (tmp4447 & tmp4448) | (tmp4447 & tmp4449) | (tmp4448 & tmp4449);
  wire tmp4451;
  assign tmp4451 = (tmp4442 & tmp4446) | (tmp4442 & tmp4450) | (tmp4446 & tmp4450);
  wire tmp4452;
  assign tmp4452 = (tmp4425 & tmp4438) | (tmp4425 & tmp4451) | (tmp4438 & tmp4451);
  wire tmp4453;
  assign tmp4453 = 1'b0;
  wire tmp4454;
  assign tmp4454 = 1'b0;
  wire tmp4455;
  assign tmp4455 = 1'b0;
  wire tmp4456;
  assign tmp4456 = (tmp4453 & tmp4454) | (tmp4453 & tmp4455) | (tmp4454 & tmp4455);
  wire tmp4457;
  assign tmp4457 = 1'b0;
  wire tmp4458;
  assign tmp4458 = 1'b1;
  wire tmp4459;
  assign tmp4459 = 1'b0;
  wire tmp4460;
  assign tmp4460 = (tmp4457 & tmp4458) | (tmp4457 & tmp4459) | (tmp4458 & tmp4459);
  wire tmp4461;
  assign tmp4461 = 1'b0;
  wire tmp4462;
  assign tmp4462 = 1'b0;
  wire tmp4463;
  assign tmp4463 = 1'b0;
  wire tmp4464;
  assign tmp4464 = (tmp4461 & tmp4462) | (tmp4461 & tmp4463) | (tmp4462 & tmp4463);
  wire tmp4465;
  assign tmp4465 = (tmp4456 & tmp4460) | (tmp4456 & tmp4464) | (tmp4460 & tmp4464);
  wire tmp4466;
  assign tmp4466 = 1'b0;
  wire tmp4467;
  assign tmp4467 = 1'b1;
  wire tmp4468;
  assign tmp4468 = 1'b0;
  wire tmp4469;
  assign tmp4469 = (tmp4466 & tmp4467) | (tmp4466 & tmp4468) | (tmp4467 & tmp4468);
  wire tmp4470;
  assign tmp4470 = 1'b1;
  wire tmp4471;
  assign tmp4471 = 1'b1;
  wire tmp4472;
  assign tmp4472 = 1'b1;
  wire tmp4473;
  assign tmp4473 = (tmp4470 & tmp4471) | (tmp4470 & tmp4472) | (tmp4471 & tmp4472);
  wire tmp4474;
  assign tmp4474 = 1'b0;
  wire tmp4475;
  assign tmp4475 = 1'b1;
  wire tmp4476;
  assign tmp4476 = 1'b0;
  wire tmp4477;
  assign tmp4477 = (tmp4474 & tmp4475) | (tmp4474 & tmp4476) | (tmp4475 & tmp4476);
  wire tmp4478;
  assign tmp4478 = (tmp4469 & tmp4473) | (tmp4469 & tmp4477) | (tmp4473 & tmp4477);
  wire tmp4479;
  assign tmp4479 = 1'b0;
  wire tmp4480;
  assign tmp4480 = 1'b0;
  wire tmp4481;
  assign tmp4481 = 1'b0;
  wire tmp4482;
  assign tmp4482 = (tmp4479 & tmp4480) | (tmp4479 & tmp4481) | (tmp4480 & tmp4481);
  wire tmp4483;
  assign tmp4483 = 1'b0;
  wire tmp4484;
  assign tmp4484 = 1'b1;
  wire tmp4485;
  assign tmp4485 = 1'b0;
  wire tmp4486;
  assign tmp4486 = (tmp4483 & tmp4484) | (tmp4483 & tmp4485) | (tmp4484 & tmp4485);
  wire tmp4487;
  assign tmp4487 = 1'b0;
  wire tmp4488;
  assign tmp4488 = 1'b0;
  wire tmp4489;
  assign tmp4489 = 1'b0;
  wire tmp4490;
  assign tmp4490 = (tmp4487 & tmp4488) | (tmp4487 & tmp4489) | (tmp4488 & tmp4489);
  wire tmp4491;
  assign tmp4491 = (tmp4482 & tmp4486) | (tmp4482 & tmp4490) | (tmp4486 & tmp4490);
  wire tmp4492;
  assign tmp4492 = (tmp4465 & tmp4478) | (tmp4465 & tmp4491) | (tmp4478 & tmp4491);
  wire tmp4493;
  assign tmp4493 = (tmp4412 & tmp4452) | (tmp4412 & tmp4492) | (tmp4452 & tmp4492);
  wire tmp4494;
  assign tmp4494 = pi3;
  wire tmp4495;
  assign tmp4495 = 1'b1;
  wire tmp4496;
  assign tmp4496 = 1'b0;
  wire tmp4497;
  assign tmp4497 = (tmp4494 & tmp4495) | (tmp4494 & tmp4496) | (tmp4495 & tmp4496);
  wire tmp4498;
  assign tmp4498 = 1'b1;
  wire tmp4499;
  assign tmp4499 = 1'b1;
  wire tmp4500;
  assign tmp4500 = 1'b1;
  wire tmp4501;
  assign tmp4501 = (tmp4498 & tmp4499) | (tmp4498 & tmp4500) | (tmp4499 & tmp4500);
  wire tmp4502;
  assign tmp4502 = 1'b0;
  wire tmp4503;
  assign tmp4503 = 1'b1;
  wire tmp4504;
  assign tmp4504 = 1'b0;
  wire tmp4505;
  assign tmp4505 = (tmp4502 & tmp4503) | (tmp4502 & tmp4504) | (tmp4503 & tmp4504);
  wire tmp4506;
  assign tmp4506 = (tmp4497 & tmp4501) | (tmp4497 & tmp4505) | (tmp4501 & tmp4505);
  wire tmp4507;
  assign tmp4507 = 1'b1;
  wire tmp4508;
  assign tmp4508 = 1'b1;
  wire tmp4509;
  assign tmp4509 = 1'b1;
  wire tmp4510;
  assign tmp4510 = (tmp4507 & tmp4508) | (tmp4507 & tmp4509) | (tmp4508 & tmp4509);
  wire tmp4511;
  assign tmp4511 = 1'b1;
  wire tmp4512;
  assign tmp4512 = 1'b1;
  wire tmp4513;
  assign tmp4513 = 1'b1;
  wire tmp4514;
  assign tmp4514 = (tmp4511 & tmp4512) | (tmp4511 & tmp4513) | (tmp4512 & tmp4513);
  wire tmp4515;
  assign tmp4515 = 1'b1;
  wire tmp4516;
  assign tmp4516 = 1'b1;
  wire tmp4517;
  assign tmp4517 = 1'b1;
  wire tmp4518;
  assign tmp4518 = (tmp4515 & tmp4516) | (tmp4515 & tmp4517) | (tmp4516 & tmp4517);
  wire tmp4519;
  assign tmp4519 = (tmp4510 & tmp4514) | (tmp4510 & tmp4518) | (tmp4514 & tmp4518);
  wire tmp4520;
  assign tmp4520 = 1'b0;
  wire tmp4521;
  assign tmp4521 = 1'b1;
  wire tmp4522;
  assign tmp4522 = 1'b0;
  wire tmp4523;
  assign tmp4523 = (tmp4520 & tmp4521) | (tmp4520 & tmp4522) | (tmp4521 & tmp4522);
  wire tmp4524;
  assign tmp4524 = 1'b1;
  wire tmp4525;
  assign tmp4525 = 1'b1;
  wire tmp4526;
  assign tmp4526 = 1'b1;
  wire tmp4527;
  assign tmp4527 = (tmp4524 & tmp4525) | (tmp4524 & tmp4526) | (tmp4525 & tmp4526);
  wire tmp4528;
  assign tmp4528 = 1'b0;
  wire tmp4529;
  assign tmp4529 = 1'b1;
  wire tmp4530;
  assign tmp4530 = 1'b0;
  wire tmp4531;
  assign tmp4531 = (tmp4528 & tmp4529) | (tmp4528 & tmp4530) | (tmp4529 & tmp4530);
  wire tmp4532;
  assign tmp4532 = (tmp4523 & tmp4527) | (tmp4523 & tmp4531) | (tmp4527 & tmp4531);
  wire tmp4533;
  assign tmp4533 = (tmp4506 & tmp4519) | (tmp4506 & tmp4532) | (tmp4519 & tmp4532);
  wire tmp4534;
  assign tmp4534 = 1'b1;
  wire tmp4535;
  assign tmp4535 = 1'b1;
  wire tmp4536;
  assign tmp4536 = 1'b1;
  wire tmp4537;
  assign tmp4537 = (tmp4534 & tmp4535) | (tmp4534 & tmp4536) | (tmp4535 & tmp4536);
  wire tmp4538;
  assign tmp4538 = 1'b1;
  wire tmp4539;
  assign tmp4539 = 1'b1;
  wire tmp4540;
  assign tmp4540 = 1'b1;
  wire tmp4541;
  assign tmp4541 = (tmp4538 & tmp4539) | (tmp4538 & tmp4540) | (tmp4539 & tmp4540);
  wire tmp4542;
  assign tmp4542 = 1'b1;
  wire tmp4543;
  assign tmp4543 = 1'b1;
  wire tmp4544;
  assign tmp4544 = 1'b1;
  wire tmp4545;
  assign tmp4545 = (tmp4542 & tmp4543) | (tmp4542 & tmp4544) | (tmp4543 & tmp4544);
  wire tmp4546;
  assign tmp4546 = (tmp4537 & tmp4541) | (tmp4537 & tmp4545) | (tmp4541 & tmp4545);
  wire tmp4547;
  assign tmp4547 = 1'b1;
  wire tmp4548;
  assign tmp4548 = 1'b1;
  wire tmp4549;
  assign tmp4549 = 1'b1;
  wire tmp4550;
  assign tmp4550 = (tmp4547 & tmp4548) | (tmp4547 & tmp4549) | (tmp4548 & tmp4549);
  wire tmp4551;
  assign tmp4551 = 1'b1;
  wire tmp4552;
  assign tmp4552 = ~pi4;
  wire tmp4553;
  assign tmp4553 = ~pi5;
  wire tmp4554;
  assign tmp4554 = (tmp4551 & tmp4552) | (tmp4551 & tmp4553) | (tmp4552 & tmp4553);
  wire tmp4555;
  assign tmp4555 = 1'b1;
  wire tmp4556;
  assign tmp4556 = ~pi5;
  wire tmp4557;
  assign tmp4557 = ~pi6;
  wire tmp4558;
  assign tmp4558 = (tmp4555 & tmp4556) | (tmp4555 & tmp4557) | (tmp4556 & tmp4557);
  wire tmp4559;
  assign tmp4559 = (tmp4550 & tmp4554) | (tmp4550 & tmp4558) | (tmp4554 & tmp4558);
  wire tmp4560;
  assign tmp4560 = 1'b1;
  wire tmp4561;
  assign tmp4561 = 1'b1;
  wire tmp4562;
  assign tmp4562 = 1'b1;
  wire tmp4563;
  assign tmp4563 = (tmp4560 & tmp4561) | (tmp4560 & tmp4562) | (tmp4561 & tmp4562);
  wire tmp4564;
  assign tmp4564 = 1'b1;
  wire tmp4565;
  assign tmp4565 = ~pi5;
  wire tmp4566;
  assign tmp4566 = ~pi6;
  wire tmp4567;
  assign tmp4567 = (tmp4564 & tmp4565) | (tmp4564 & tmp4566) | (tmp4565 & tmp4566);
  wire tmp4568;
  assign tmp4568 = 1'b1;
  wire tmp4569;
  assign tmp4569 = ~pi6;
  wire tmp4570;
  assign tmp4570 = ~pi7;
  wire tmp4571;
  assign tmp4571 = (tmp4568 & tmp4569) | (tmp4568 & tmp4570) | (tmp4569 & tmp4570);
  wire tmp4572;
  assign tmp4572 = (tmp4563 & tmp4567) | (tmp4563 & tmp4571) | (tmp4567 & tmp4571);
  wire tmp4573;
  assign tmp4573 = (tmp4546 & tmp4559) | (tmp4546 & tmp4572) | (tmp4559 & tmp4572);
  wire tmp4574;
  assign tmp4574 = 1'b0;
  wire tmp4575;
  assign tmp4575 = 1'b1;
  wire tmp4576;
  assign tmp4576 = 1'b0;
  wire tmp4577;
  assign tmp4577 = (tmp4574 & tmp4575) | (tmp4574 & tmp4576) | (tmp4575 & tmp4576);
  wire tmp4578;
  assign tmp4578 = 1'b1;
  wire tmp4579;
  assign tmp4579 = 1'b1;
  wire tmp4580;
  assign tmp4580 = 1'b1;
  wire tmp4581;
  assign tmp4581 = (tmp4578 & tmp4579) | (tmp4578 & tmp4580) | (tmp4579 & tmp4580);
  wire tmp4582;
  assign tmp4582 = 1'b0;
  wire tmp4583;
  assign tmp4583 = 1'b1;
  wire tmp4584;
  assign tmp4584 = 1'b0;
  wire tmp4585;
  assign tmp4585 = (tmp4582 & tmp4583) | (tmp4582 & tmp4584) | (tmp4583 & tmp4584);
  wire tmp4586;
  assign tmp4586 = (tmp4577 & tmp4581) | (tmp4577 & tmp4585) | (tmp4581 & tmp4585);
  wire tmp4587;
  assign tmp4587 = 1'b1;
  wire tmp4588;
  assign tmp4588 = 1'b1;
  wire tmp4589;
  assign tmp4589 = 1'b1;
  wire tmp4590;
  assign tmp4590 = (tmp4587 & tmp4588) | (tmp4587 & tmp4589) | (tmp4588 & tmp4589);
  wire tmp4591;
  assign tmp4591 = 1'b1;
  wire tmp4592;
  assign tmp4592 = ~pi5;
  wire tmp4593;
  assign tmp4593 = ~pi6;
  wire tmp4594;
  assign tmp4594 = (tmp4591 & tmp4592) | (tmp4591 & tmp4593) | (tmp4592 & tmp4593);
  wire tmp4595;
  assign tmp4595 = 1'b1;
  wire tmp4596;
  assign tmp4596 = ~pi6;
  wire tmp4597;
  assign tmp4597 = ~pi7;
  wire tmp4598;
  assign tmp4598 = (tmp4595 & tmp4596) | (tmp4595 & tmp4597) | (tmp4596 & tmp4597);
  wire tmp4599;
  assign tmp4599 = (tmp4590 & tmp4594) | (tmp4590 & tmp4598) | (tmp4594 & tmp4598);
  wire tmp4600;
  assign tmp4600 = 1'b0;
  wire tmp4601;
  assign tmp4601 = 1'b1;
  wire tmp4602;
  assign tmp4602 = 1'b0;
  wire tmp4603;
  assign tmp4603 = (tmp4600 & tmp4601) | (tmp4600 & tmp4602) | (tmp4601 & tmp4602);
  wire tmp4604;
  assign tmp4604 = 1'b1;
  wire tmp4605;
  assign tmp4605 = ~pi6;
  wire tmp4606;
  assign tmp4606 = ~pi7;
  wire tmp4607;
  assign tmp4607 = (tmp4604 & tmp4605) | (tmp4604 & tmp4606) | (tmp4605 & tmp4606);
  wire tmp4608;
  assign tmp4608 = 1'b0;
  wire tmp4609;
  assign tmp4609 = ~pi7;
  wire tmp4610;
  assign tmp4610 = 1'b0;
  wire tmp4611;
  assign tmp4611 = (tmp4608 & tmp4609) | (tmp4608 & tmp4610) | (tmp4609 & tmp4610);
  wire tmp4612;
  assign tmp4612 = (tmp4603 & tmp4607) | (tmp4603 & tmp4611) | (tmp4607 & tmp4611);
  wire tmp4613;
  assign tmp4613 = (tmp4586 & tmp4599) | (tmp4586 & tmp4612) | (tmp4599 & tmp4612);
  wire tmp4614;
  assign tmp4614 = (tmp4533 & tmp4573) | (tmp4533 & tmp4613) | (tmp4573 & tmp4613);
  wire tmp4615;
  assign tmp4615 = 1'b0;
  wire tmp4616;
  assign tmp4616 = 1'b0;
  wire tmp4617;
  assign tmp4617 = 1'b0;
  wire tmp4618;
  assign tmp4618 = (tmp4615 & tmp4616) | (tmp4615 & tmp4617) | (tmp4616 & tmp4617);
  wire tmp4619;
  assign tmp4619 = 1'b0;
  wire tmp4620;
  assign tmp4620 = 1'b1;
  wire tmp4621;
  assign tmp4621 = 1'b0;
  wire tmp4622;
  assign tmp4622 = (tmp4619 & tmp4620) | (tmp4619 & tmp4621) | (tmp4620 & tmp4621);
  wire tmp4623;
  assign tmp4623 = 1'b0;
  wire tmp4624;
  assign tmp4624 = 1'b0;
  wire tmp4625;
  assign tmp4625 = 1'b0;
  wire tmp4626;
  assign tmp4626 = (tmp4623 & tmp4624) | (tmp4623 & tmp4625) | (tmp4624 & tmp4625);
  wire tmp4627;
  assign tmp4627 = (tmp4618 & tmp4622) | (tmp4618 & tmp4626) | (tmp4622 & tmp4626);
  wire tmp4628;
  assign tmp4628 = 1'b0;
  wire tmp4629;
  assign tmp4629 = 1'b1;
  wire tmp4630;
  assign tmp4630 = 1'b0;
  wire tmp4631;
  assign tmp4631 = (tmp4628 & tmp4629) | (tmp4628 & tmp4630) | (tmp4629 & tmp4630);
  wire tmp4632;
  assign tmp4632 = 1'b1;
  wire tmp4633;
  assign tmp4633 = 1'b1;
  wire tmp4634;
  assign tmp4634 = 1'b1;
  wire tmp4635;
  assign tmp4635 = (tmp4632 & tmp4633) | (tmp4632 & tmp4634) | (tmp4633 & tmp4634);
  wire tmp4636;
  assign tmp4636 = 1'b0;
  wire tmp4637;
  assign tmp4637 = 1'b1;
  wire tmp4638;
  assign tmp4638 = 1'b0;
  wire tmp4639;
  assign tmp4639 = (tmp4636 & tmp4637) | (tmp4636 & tmp4638) | (tmp4637 & tmp4638);
  wire tmp4640;
  assign tmp4640 = (tmp4631 & tmp4635) | (tmp4631 & tmp4639) | (tmp4635 & tmp4639);
  wire tmp4641;
  assign tmp4641 = 1'b0;
  wire tmp4642;
  assign tmp4642 = 1'b0;
  wire tmp4643;
  assign tmp4643 = 1'b0;
  wire tmp4644;
  assign tmp4644 = (tmp4641 & tmp4642) | (tmp4641 & tmp4643) | (tmp4642 & tmp4643);
  wire tmp4645;
  assign tmp4645 = 1'b0;
  wire tmp4646;
  assign tmp4646 = 1'b1;
  wire tmp4647;
  assign tmp4647 = 1'b0;
  wire tmp4648;
  assign tmp4648 = (tmp4645 & tmp4646) | (tmp4645 & tmp4647) | (tmp4646 & tmp4647);
  wire tmp4649;
  assign tmp4649 = 1'b0;
  wire tmp4650;
  assign tmp4650 = 1'b0;
  wire tmp4651;
  assign tmp4651 = 1'b0;
  wire tmp4652;
  assign tmp4652 = (tmp4649 & tmp4650) | (tmp4649 & tmp4651) | (tmp4650 & tmp4651);
  wire tmp4653;
  assign tmp4653 = (tmp4644 & tmp4648) | (tmp4644 & tmp4652) | (tmp4648 & tmp4652);
  wire tmp4654;
  assign tmp4654 = (tmp4627 & tmp4640) | (tmp4627 & tmp4653) | (tmp4640 & tmp4653);
  wire tmp4655;
  assign tmp4655 = 1'b0;
  wire tmp4656;
  assign tmp4656 = 1'b1;
  wire tmp4657;
  assign tmp4657 = 1'b0;
  wire tmp4658;
  assign tmp4658 = (tmp4655 & tmp4656) | (tmp4655 & tmp4657) | (tmp4656 & tmp4657);
  wire tmp4659;
  assign tmp4659 = 1'b1;
  wire tmp4660;
  assign tmp4660 = 1'b1;
  wire tmp4661;
  assign tmp4661 = 1'b1;
  wire tmp4662;
  assign tmp4662 = (tmp4659 & tmp4660) | (tmp4659 & tmp4661) | (tmp4660 & tmp4661);
  wire tmp4663;
  assign tmp4663 = 1'b0;
  wire tmp4664;
  assign tmp4664 = 1'b1;
  wire tmp4665;
  assign tmp4665 = 1'b0;
  wire tmp4666;
  assign tmp4666 = (tmp4663 & tmp4664) | (tmp4663 & tmp4665) | (tmp4664 & tmp4665);
  wire tmp4667;
  assign tmp4667 = (tmp4658 & tmp4662) | (tmp4658 & tmp4666) | (tmp4662 & tmp4666);
  wire tmp4668;
  assign tmp4668 = 1'b1;
  wire tmp4669;
  assign tmp4669 = 1'b1;
  wire tmp4670;
  assign tmp4670 = 1'b1;
  wire tmp4671;
  assign tmp4671 = (tmp4668 & tmp4669) | (tmp4668 & tmp4670) | (tmp4669 & tmp4670);
  wire tmp4672;
  assign tmp4672 = 1'b1;
  wire tmp4673;
  assign tmp4673 = ~pi5;
  wire tmp4674;
  assign tmp4674 = ~pi6;
  wire tmp4675;
  assign tmp4675 = (tmp4672 & tmp4673) | (tmp4672 & tmp4674) | (tmp4673 & tmp4674);
  wire tmp4676;
  assign tmp4676 = 1'b1;
  wire tmp4677;
  assign tmp4677 = ~pi6;
  wire tmp4678;
  assign tmp4678 = ~pi7;
  wire tmp4679;
  assign tmp4679 = (tmp4676 & tmp4677) | (tmp4676 & tmp4678) | (tmp4677 & tmp4678);
  wire tmp4680;
  assign tmp4680 = (tmp4671 & tmp4675) | (tmp4671 & tmp4679) | (tmp4675 & tmp4679);
  wire tmp4681;
  assign tmp4681 = 1'b0;
  wire tmp4682;
  assign tmp4682 = 1'b1;
  wire tmp4683;
  assign tmp4683 = 1'b0;
  wire tmp4684;
  assign tmp4684 = (tmp4681 & tmp4682) | (tmp4681 & tmp4683) | (tmp4682 & tmp4683);
  wire tmp4685;
  assign tmp4685 = 1'b1;
  wire tmp4686;
  assign tmp4686 = ~pi6;
  wire tmp4687;
  assign tmp4687 = ~pi7;
  wire tmp4688;
  assign tmp4688 = (tmp4685 & tmp4686) | (tmp4685 & tmp4687) | (tmp4686 & tmp4687);
  wire tmp4689;
  assign tmp4689 = 1'b0;
  wire tmp4690;
  assign tmp4690 = ~pi7;
  wire tmp4691;
  assign tmp4691 = 1'b0;
  wire tmp4692;
  assign tmp4692 = (tmp4689 & tmp4690) | (tmp4689 & tmp4691) | (tmp4690 & tmp4691);
  wire tmp4693;
  assign tmp4693 = (tmp4684 & tmp4688) | (tmp4684 & tmp4692) | (tmp4688 & tmp4692);
  wire tmp4694;
  assign tmp4694 = (tmp4667 & tmp4680) | (tmp4667 & tmp4693) | (tmp4680 & tmp4693);
  wire tmp4695;
  assign tmp4695 = 1'b0;
  wire tmp4696;
  assign tmp4696 = 1'b0;
  wire tmp4697;
  assign tmp4697 = 1'b0;
  wire tmp4698;
  assign tmp4698 = (tmp4695 & tmp4696) | (tmp4695 & tmp4697) | (tmp4696 & tmp4697);
  wire tmp4699;
  assign tmp4699 = 1'b0;
  wire tmp4700;
  assign tmp4700 = 1'b1;
  wire tmp4701;
  assign tmp4701 = 1'b0;
  wire tmp4702;
  assign tmp4702 = (tmp4699 & tmp4700) | (tmp4699 & tmp4701) | (tmp4700 & tmp4701);
  wire tmp4703;
  assign tmp4703 = 1'b0;
  wire tmp4704;
  assign tmp4704 = 1'b0;
  wire tmp4705;
  assign tmp4705 = 1'b0;
  wire tmp4706;
  assign tmp4706 = (tmp4703 & tmp4704) | (tmp4703 & tmp4705) | (tmp4704 & tmp4705);
  wire tmp4707;
  assign tmp4707 = (tmp4698 & tmp4702) | (tmp4698 & tmp4706) | (tmp4702 & tmp4706);
  wire tmp4708;
  assign tmp4708 = 1'b0;
  wire tmp4709;
  assign tmp4709 = 1'b1;
  wire tmp4710;
  assign tmp4710 = 1'b0;
  wire tmp4711;
  assign tmp4711 = (tmp4708 & tmp4709) | (tmp4708 & tmp4710) | (tmp4709 & tmp4710);
  wire tmp4712;
  assign tmp4712 = 1'b1;
  wire tmp4713;
  assign tmp4713 = ~pi6;
  wire tmp4714;
  assign tmp4714 = ~pi7;
  wire tmp4715;
  assign tmp4715 = (tmp4712 & tmp4713) | (tmp4712 & tmp4714) | (tmp4713 & tmp4714);
  wire tmp4716;
  assign tmp4716 = 1'b0;
  wire tmp4717;
  assign tmp4717 = ~pi7;
  wire tmp4718;
  assign tmp4718 = 1'b0;
  wire tmp4719;
  assign tmp4719 = (tmp4716 & tmp4717) | (tmp4716 & tmp4718) | (tmp4717 & tmp4718);
  wire tmp4720;
  assign tmp4720 = (tmp4711 & tmp4715) | (tmp4711 & tmp4719) | (tmp4715 & tmp4719);
  wire tmp4721;
  assign tmp4721 = 1'b0;
  wire tmp4722;
  assign tmp4722 = 1'b0;
  wire tmp4723;
  assign tmp4723 = 1'b0;
  wire tmp4724;
  assign tmp4724 = (tmp4721 & tmp4722) | (tmp4721 & tmp4723) | (tmp4722 & tmp4723);
  wire tmp4725;
  assign tmp4725 = 1'b0;
  wire tmp4726;
  assign tmp4726 = ~pi7;
  wire tmp4727;
  assign tmp4727 = 1'b0;
  wire tmp4728;
  assign tmp4728 = (tmp4725 & tmp4726) | (tmp4725 & tmp4727) | (tmp4726 & tmp4727);
  wire tmp4729;
  assign tmp4729 = 1'b0;
  wire tmp4730;
  assign tmp4730 = 1'b0;
  wire tmp4731;
  assign tmp4731 = 1'b0;
  wire tmp4732;
  assign tmp4732 = (tmp4729 & tmp4730) | (tmp4729 & tmp4731) | (tmp4730 & tmp4731);
  wire tmp4733;
  assign tmp4733 = (tmp4724 & tmp4728) | (tmp4724 & tmp4732) | (tmp4728 & tmp4732);
  wire tmp4734;
  assign tmp4734 = (tmp4707 & tmp4720) | (tmp4707 & tmp4733) | (tmp4720 & tmp4733);
  wire tmp4735;
  assign tmp4735 = (tmp4654 & tmp4694) | (tmp4654 & tmp4734) | (tmp4694 & tmp4734);
  wire tmp4736;
  assign tmp4736 = (tmp4493 & tmp4614) | (tmp4493 & tmp4735) | (tmp4614 & tmp4735);
  wire tmp4737;
  assign tmp4737 = pi3;
  wire tmp4738;
  assign tmp4738 = 1'b1;
  wire tmp4739;
  assign tmp4739 = 1'b0;
  wire tmp4740;
  assign tmp4740 = (tmp4737 & tmp4738) | (tmp4737 & tmp4739) | (tmp4738 & tmp4739);
  wire tmp4741;
  assign tmp4741 = 1'b1;
  wire tmp4742;
  assign tmp4742 = 1'b1;
  wire tmp4743;
  assign tmp4743 = 1'b1;
  wire tmp4744;
  assign tmp4744 = (tmp4741 & tmp4742) | (tmp4741 & tmp4743) | (tmp4742 & tmp4743);
  wire tmp4745;
  assign tmp4745 = 1'b0;
  wire tmp4746;
  assign tmp4746 = 1'b1;
  wire tmp4747;
  assign tmp4747 = 1'b0;
  wire tmp4748;
  assign tmp4748 = (tmp4745 & tmp4746) | (tmp4745 & tmp4747) | (tmp4746 & tmp4747);
  wire tmp4749;
  assign tmp4749 = (tmp4740 & tmp4744) | (tmp4740 & tmp4748) | (tmp4744 & tmp4748);
  wire tmp4750;
  assign tmp4750 = 1'b1;
  wire tmp4751;
  assign tmp4751 = 1'b1;
  wire tmp4752;
  assign tmp4752 = 1'b1;
  wire tmp4753;
  assign tmp4753 = (tmp4750 & tmp4751) | (tmp4750 & tmp4752) | (tmp4751 & tmp4752);
  wire tmp4754;
  assign tmp4754 = 1'b1;
  wire tmp4755;
  assign tmp4755 = 1'b1;
  wire tmp4756;
  assign tmp4756 = 1'b1;
  wire tmp4757;
  assign tmp4757 = (tmp4754 & tmp4755) | (tmp4754 & tmp4756) | (tmp4755 & tmp4756);
  wire tmp4758;
  assign tmp4758 = 1'b1;
  wire tmp4759;
  assign tmp4759 = 1'b1;
  wire tmp4760;
  assign tmp4760 = 1'b1;
  wire tmp4761;
  assign tmp4761 = (tmp4758 & tmp4759) | (tmp4758 & tmp4760) | (tmp4759 & tmp4760);
  wire tmp4762;
  assign tmp4762 = (tmp4753 & tmp4757) | (tmp4753 & tmp4761) | (tmp4757 & tmp4761);
  wire tmp4763;
  assign tmp4763 = 1'b0;
  wire tmp4764;
  assign tmp4764 = 1'b1;
  wire tmp4765;
  assign tmp4765 = 1'b0;
  wire tmp4766;
  assign tmp4766 = (tmp4763 & tmp4764) | (tmp4763 & tmp4765) | (tmp4764 & tmp4765);
  wire tmp4767;
  assign tmp4767 = 1'b1;
  wire tmp4768;
  assign tmp4768 = 1'b1;
  wire tmp4769;
  assign tmp4769 = 1'b1;
  wire tmp4770;
  assign tmp4770 = (tmp4767 & tmp4768) | (tmp4767 & tmp4769) | (tmp4768 & tmp4769);
  wire tmp4771;
  assign tmp4771 = 1'b0;
  wire tmp4772;
  assign tmp4772 = 1'b1;
  wire tmp4773;
  assign tmp4773 = 1'b0;
  wire tmp4774;
  assign tmp4774 = (tmp4771 & tmp4772) | (tmp4771 & tmp4773) | (tmp4772 & tmp4773);
  wire tmp4775;
  assign tmp4775 = (tmp4766 & tmp4770) | (tmp4766 & tmp4774) | (tmp4770 & tmp4774);
  wire tmp4776;
  assign tmp4776 = (tmp4749 & tmp4762) | (tmp4749 & tmp4775) | (tmp4762 & tmp4775);
  wire tmp4777;
  assign tmp4777 = 1'b1;
  wire tmp4778;
  assign tmp4778 = 1'b1;
  wire tmp4779;
  assign tmp4779 = 1'b1;
  wire tmp4780;
  assign tmp4780 = (tmp4777 & tmp4778) | (tmp4777 & tmp4779) | (tmp4778 & tmp4779);
  wire tmp4781;
  assign tmp4781 = 1'b1;
  wire tmp4782;
  assign tmp4782 = 1'b1;
  wire tmp4783;
  assign tmp4783 = 1'b1;
  wire tmp4784;
  assign tmp4784 = (tmp4781 & tmp4782) | (tmp4781 & tmp4783) | (tmp4782 & tmp4783);
  wire tmp4785;
  assign tmp4785 = 1'b1;
  wire tmp4786;
  assign tmp4786 = 1'b1;
  wire tmp4787;
  assign tmp4787 = 1'b1;
  wire tmp4788;
  assign tmp4788 = (tmp4785 & tmp4786) | (tmp4785 & tmp4787) | (tmp4786 & tmp4787);
  wire tmp4789;
  assign tmp4789 = (tmp4780 & tmp4784) | (tmp4780 & tmp4788) | (tmp4784 & tmp4788);
  wire tmp4790;
  assign tmp4790 = 1'b1;
  wire tmp4791;
  assign tmp4791 = 1'b1;
  wire tmp4792;
  assign tmp4792 = 1'b1;
  wire tmp4793;
  assign tmp4793 = (tmp4790 & tmp4791) | (tmp4790 & tmp4792) | (tmp4791 & tmp4792);
  wire tmp4794;
  assign tmp4794 = 1'b1;
  wire tmp4795;
  assign tmp4795 = ~pi4;
  wire tmp4796;
  assign tmp4796 = ~pi5;
  wire tmp4797;
  assign tmp4797 = (tmp4794 & tmp4795) | (tmp4794 & tmp4796) | (tmp4795 & tmp4796);
  wire tmp4798;
  assign tmp4798 = 1'b1;
  wire tmp4799;
  assign tmp4799 = ~pi5;
  wire tmp4800;
  assign tmp4800 = ~pi6;
  wire tmp4801;
  assign tmp4801 = (tmp4798 & tmp4799) | (tmp4798 & tmp4800) | (tmp4799 & tmp4800);
  wire tmp4802;
  assign tmp4802 = (tmp4793 & tmp4797) | (tmp4793 & tmp4801) | (tmp4797 & tmp4801);
  wire tmp4803;
  assign tmp4803 = 1'b1;
  wire tmp4804;
  assign tmp4804 = 1'b1;
  wire tmp4805;
  assign tmp4805 = 1'b1;
  wire tmp4806;
  assign tmp4806 = (tmp4803 & tmp4804) | (tmp4803 & tmp4805) | (tmp4804 & tmp4805);
  wire tmp4807;
  assign tmp4807 = 1'b1;
  wire tmp4808;
  assign tmp4808 = ~pi5;
  wire tmp4809;
  assign tmp4809 = ~pi6;
  wire tmp4810;
  assign tmp4810 = (tmp4807 & tmp4808) | (tmp4807 & tmp4809) | (tmp4808 & tmp4809);
  wire tmp4811;
  assign tmp4811 = 1'b1;
  wire tmp4812;
  assign tmp4812 = ~pi6;
  wire tmp4813;
  assign tmp4813 = ~pi7;
  wire tmp4814;
  assign tmp4814 = (tmp4811 & tmp4812) | (tmp4811 & tmp4813) | (tmp4812 & tmp4813);
  wire tmp4815;
  assign tmp4815 = (tmp4806 & tmp4810) | (tmp4806 & tmp4814) | (tmp4810 & tmp4814);
  wire tmp4816;
  assign tmp4816 = (tmp4789 & tmp4802) | (tmp4789 & tmp4815) | (tmp4802 & tmp4815);
  wire tmp4817;
  assign tmp4817 = 1'b0;
  wire tmp4818;
  assign tmp4818 = 1'b1;
  wire tmp4819;
  assign tmp4819 = 1'b0;
  wire tmp4820;
  assign tmp4820 = (tmp4817 & tmp4818) | (tmp4817 & tmp4819) | (tmp4818 & tmp4819);
  wire tmp4821;
  assign tmp4821 = 1'b1;
  wire tmp4822;
  assign tmp4822 = 1'b1;
  wire tmp4823;
  assign tmp4823 = 1'b1;
  wire tmp4824;
  assign tmp4824 = (tmp4821 & tmp4822) | (tmp4821 & tmp4823) | (tmp4822 & tmp4823);
  wire tmp4825;
  assign tmp4825 = 1'b0;
  wire tmp4826;
  assign tmp4826 = 1'b1;
  wire tmp4827;
  assign tmp4827 = 1'b0;
  wire tmp4828;
  assign tmp4828 = (tmp4825 & tmp4826) | (tmp4825 & tmp4827) | (tmp4826 & tmp4827);
  wire tmp4829;
  assign tmp4829 = (tmp4820 & tmp4824) | (tmp4820 & tmp4828) | (tmp4824 & tmp4828);
  wire tmp4830;
  assign tmp4830 = 1'b1;
  wire tmp4831;
  assign tmp4831 = 1'b1;
  wire tmp4832;
  assign tmp4832 = 1'b1;
  wire tmp4833;
  assign tmp4833 = (tmp4830 & tmp4831) | (tmp4830 & tmp4832) | (tmp4831 & tmp4832);
  wire tmp4834;
  assign tmp4834 = 1'b1;
  wire tmp4835;
  assign tmp4835 = ~pi5;
  wire tmp4836;
  assign tmp4836 = ~pi6;
  wire tmp4837;
  assign tmp4837 = (tmp4834 & tmp4835) | (tmp4834 & tmp4836) | (tmp4835 & tmp4836);
  wire tmp4838;
  assign tmp4838 = 1'b1;
  wire tmp4839;
  assign tmp4839 = ~pi6;
  wire tmp4840;
  assign tmp4840 = ~pi7;
  wire tmp4841;
  assign tmp4841 = (tmp4838 & tmp4839) | (tmp4838 & tmp4840) | (tmp4839 & tmp4840);
  wire tmp4842;
  assign tmp4842 = (tmp4833 & tmp4837) | (tmp4833 & tmp4841) | (tmp4837 & tmp4841);
  wire tmp4843;
  assign tmp4843 = 1'b0;
  wire tmp4844;
  assign tmp4844 = 1'b1;
  wire tmp4845;
  assign tmp4845 = 1'b0;
  wire tmp4846;
  assign tmp4846 = (tmp4843 & tmp4844) | (tmp4843 & tmp4845) | (tmp4844 & tmp4845);
  wire tmp4847;
  assign tmp4847 = 1'b1;
  wire tmp4848;
  assign tmp4848 = ~pi6;
  wire tmp4849;
  assign tmp4849 = ~pi7;
  wire tmp4850;
  assign tmp4850 = (tmp4847 & tmp4848) | (tmp4847 & tmp4849) | (tmp4848 & tmp4849);
  wire tmp4851;
  assign tmp4851 = 1'b0;
  wire tmp4852;
  assign tmp4852 = ~pi7;
  wire tmp4853;
  assign tmp4853 = 1'b0;
  wire tmp4854;
  assign tmp4854 = (tmp4851 & tmp4852) | (tmp4851 & tmp4853) | (tmp4852 & tmp4853);
  wire tmp4855;
  assign tmp4855 = (tmp4846 & tmp4850) | (tmp4846 & tmp4854) | (tmp4850 & tmp4854);
  wire tmp4856;
  assign tmp4856 = (tmp4829 & tmp4842) | (tmp4829 & tmp4855) | (tmp4842 & tmp4855);
  wire tmp4857;
  assign tmp4857 = (tmp4776 & tmp4816) | (tmp4776 & tmp4856) | (tmp4816 & tmp4856);
  wire tmp4858;
  assign tmp4858 = 1'b1;
  wire tmp4859;
  assign tmp4859 = 1'b1;
  wire tmp4860;
  assign tmp4860 = 1'b1;
  wire tmp4861;
  assign tmp4861 = (tmp4858 & tmp4859) | (tmp4858 & tmp4860) | (tmp4859 & tmp4860);
  wire tmp4862;
  assign tmp4862 = 1'b1;
  wire tmp4863;
  assign tmp4863 = 1'b1;
  wire tmp4864;
  assign tmp4864 = 1'b1;
  wire tmp4865;
  assign tmp4865 = (tmp4862 & tmp4863) | (tmp4862 & tmp4864) | (tmp4863 & tmp4864);
  wire tmp4866;
  assign tmp4866 = 1'b1;
  wire tmp4867;
  assign tmp4867 = 1'b1;
  wire tmp4868;
  assign tmp4868 = 1'b1;
  wire tmp4869;
  assign tmp4869 = (tmp4866 & tmp4867) | (tmp4866 & tmp4868) | (tmp4867 & tmp4868);
  wire tmp4870;
  assign tmp4870 = (tmp4861 & tmp4865) | (tmp4861 & tmp4869) | (tmp4865 & tmp4869);
  wire tmp4871;
  assign tmp4871 = 1'b1;
  wire tmp4872;
  assign tmp4872 = 1'b1;
  wire tmp4873;
  assign tmp4873 = 1'b1;
  wire tmp4874;
  assign tmp4874 = (tmp4871 & tmp4872) | (tmp4871 & tmp4873) | (tmp4872 & tmp4873);
  wire tmp4875;
  assign tmp4875 = 1'b1;
  wire tmp4876;
  assign tmp4876 = ~pi4;
  wire tmp4877;
  assign tmp4877 = ~pi5;
  wire tmp4878;
  assign tmp4878 = (tmp4875 & tmp4876) | (tmp4875 & tmp4877) | (tmp4876 & tmp4877);
  wire tmp4879;
  assign tmp4879 = 1'b1;
  wire tmp4880;
  assign tmp4880 = ~pi5;
  wire tmp4881;
  assign tmp4881 = ~pi6;
  wire tmp4882;
  assign tmp4882 = (tmp4879 & tmp4880) | (tmp4879 & tmp4881) | (tmp4880 & tmp4881);
  wire tmp4883;
  assign tmp4883 = (tmp4874 & tmp4878) | (tmp4874 & tmp4882) | (tmp4878 & tmp4882);
  wire tmp4884;
  assign tmp4884 = 1'b1;
  wire tmp4885;
  assign tmp4885 = 1'b1;
  wire tmp4886;
  assign tmp4886 = 1'b1;
  wire tmp4887;
  assign tmp4887 = (tmp4884 & tmp4885) | (tmp4884 & tmp4886) | (tmp4885 & tmp4886);
  wire tmp4888;
  assign tmp4888 = 1'b1;
  wire tmp4889;
  assign tmp4889 = ~pi5;
  wire tmp4890;
  assign tmp4890 = ~pi6;
  wire tmp4891;
  assign tmp4891 = (tmp4888 & tmp4889) | (tmp4888 & tmp4890) | (tmp4889 & tmp4890);
  wire tmp4892;
  assign tmp4892 = 1'b1;
  wire tmp4893;
  assign tmp4893 = ~pi6;
  wire tmp4894;
  assign tmp4894 = ~pi7;
  wire tmp4895;
  assign tmp4895 = (tmp4892 & tmp4893) | (tmp4892 & tmp4894) | (tmp4893 & tmp4894);
  wire tmp4896;
  assign tmp4896 = (tmp4887 & tmp4891) | (tmp4887 & tmp4895) | (tmp4891 & tmp4895);
  wire tmp4897;
  assign tmp4897 = (tmp4870 & tmp4883) | (tmp4870 & tmp4896) | (tmp4883 & tmp4896);
  wire tmp4898;
  assign tmp4898 = 1'b1;
  wire tmp4899;
  assign tmp4899 = 1'b1;
  wire tmp4900;
  assign tmp4900 = 1'b1;
  wire tmp4901;
  assign tmp4901 = (tmp4898 & tmp4899) | (tmp4898 & tmp4900) | (tmp4899 & tmp4900);
  wire tmp4902;
  assign tmp4902 = 1'b1;
  wire tmp4903;
  assign tmp4903 = ~pi4;
  wire tmp4904;
  assign tmp4904 = ~pi5;
  wire tmp4905;
  assign tmp4905 = (tmp4902 & tmp4903) | (tmp4902 & tmp4904) | (tmp4903 & tmp4904);
  wire tmp4906;
  assign tmp4906 = 1'b1;
  wire tmp4907;
  assign tmp4907 = ~pi5;
  wire tmp4908;
  assign tmp4908 = ~pi6;
  wire tmp4909;
  assign tmp4909 = (tmp4906 & tmp4907) | (tmp4906 & tmp4908) | (tmp4907 & tmp4908);
  wire tmp4910;
  assign tmp4910 = (tmp4901 & tmp4905) | (tmp4901 & tmp4909) | (tmp4905 & tmp4909);
  wire tmp4911;
  assign tmp4911 = 1'b1;
  wire tmp4912;
  assign tmp4912 = ~pi4;
  wire tmp4913;
  assign tmp4913 = ~pi5;
  wire tmp4914;
  assign tmp4914 = (tmp4911 & tmp4912) | (tmp4911 & tmp4913) | (tmp4912 & tmp4913);
  wire tmp4915;
  assign tmp4915 = ~pi4;
  wire tmp4916;
  assign tmp4916 = 1'b1;
  wire tmp4917;
  assign tmp4917 = 1'b1;
  wire tmp4918;
  assign tmp4918 = (tmp4915 & tmp4916) | (tmp4915 & tmp4917) | (tmp4916 & tmp4917);
  wire tmp4919;
  assign tmp4919 = ~pi5;
  wire tmp4920;
  assign tmp4920 = 1'b1;
  wire tmp4921;
  assign tmp4921 = 1'b1;
  wire tmp4922;
  assign tmp4922 = (tmp4919 & tmp4920) | (tmp4919 & tmp4921) | (tmp4920 & tmp4921);
  wire tmp4923;
  assign tmp4923 = (tmp4914 & tmp4918) | (tmp4914 & tmp4922) | (tmp4918 & tmp4922);
  wire tmp4924;
  assign tmp4924 = 1'b1;
  wire tmp4925;
  assign tmp4925 = ~pi5;
  wire tmp4926;
  assign tmp4926 = ~pi6;
  wire tmp4927;
  assign tmp4927 = (tmp4924 & tmp4925) | (tmp4924 & tmp4926) | (tmp4925 & tmp4926);
  wire tmp4928;
  assign tmp4928 = ~pi5;
  wire tmp4929;
  assign tmp4929 = 1'b1;
  wire tmp4930;
  assign tmp4930 = 1'b1;
  wire tmp4931;
  assign tmp4931 = (tmp4928 & tmp4929) | (tmp4928 & tmp4930) | (tmp4929 & tmp4930);
  wire tmp4932;
  assign tmp4932 = ~pi6;
  wire tmp4933;
  assign tmp4933 = 1'b1;
  wire tmp4934;
  assign tmp4934 = 1'b1;
  wire tmp4935;
  assign tmp4935 = (tmp4932 & tmp4933) | (tmp4932 & tmp4934) | (tmp4933 & tmp4934);
  wire tmp4936;
  assign tmp4936 = (tmp4927 & tmp4931) | (tmp4927 & tmp4935) | (tmp4931 & tmp4935);
  wire tmp4937;
  assign tmp4937 = (tmp4910 & tmp4923) | (tmp4910 & tmp4936) | (tmp4923 & tmp4936);
  wire tmp4938;
  assign tmp4938 = 1'b1;
  wire tmp4939;
  assign tmp4939 = 1'b1;
  wire tmp4940;
  assign tmp4940 = 1'b1;
  wire tmp4941;
  assign tmp4941 = (tmp4938 & tmp4939) | (tmp4938 & tmp4940) | (tmp4939 & tmp4940);
  wire tmp4942;
  assign tmp4942 = 1'b1;
  wire tmp4943;
  assign tmp4943 = ~pi5;
  wire tmp4944;
  assign tmp4944 = ~pi6;
  wire tmp4945;
  assign tmp4945 = (tmp4942 & tmp4943) | (tmp4942 & tmp4944) | (tmp4943 & tmp4944);
  wire tmp4946;
  assign tmp4946 = 1'b1;
  wire tmp4947;
  assign tmp4947 = ~pi6;
  wire tmp4948;
  assign tmp4948 = ~pi7;
  wire tmp4949;
  assign tmp4949 = (tmp4946 & tmp4947) | (tmp4946 & tmp4948) | (tmp4947 & tmp4948);
  wire tmp4950;
  assign tmp4950 = (tmp4941 & tmp4945) | (tmp4941 & tmp4949) | (tmp4945 & tmp4949);
  wire tmp4951;
  assign tmp4951 = 1'b1;
  wire tmp4952;
  assign tmp4952 = ~pi5;
  wire tmp4953;
  assign tmp4953 = ~pi6;
  wire tmp4954;
  assign tmp4954 = (tmp4951 & tmp4952) | (tmp4951 & tmp4953) | (tmp4952 & tmp4953);
  wire tmp4955;
  assign tmp4955 = ~pi5;
  wire tmp4956;
  assign tmp4956 = 1'b1;
  wire tmp4957;
  assign tmp4957 = 1'b1;
  wire tmp4958;
  assign tmp4958 = (tmp4955 & tmp4956) | (tmp4955 & tmp4957) | (tmp4956 & tmp4957);
  wire tmp4959;
  assign tmp4959 = ~pi6;
  wire tmp4960;
  assign tmp4960 = 1'b1;
  wire tmp4961;
  assign tmp4961 = 1'b1;
  wire tmp4962;
  assign tmp4962 = (tmp4959 & tmp4960) | (tmp4959 & tmp4961) | (tmp4960 & tmp4961);
  wire tmp4963;
  assign tmp4963 = (tmp4954 & tmp4958) | (tmp4954 & tmp4962) | (tmp4958 & tmp4962);
  wire tmp4964;
  assign tmp4964 = 1'b1;
  wire tmp4965;
  assign tmp4965 = ~pi6;
  wire tmp4966;
  assign tmp4966 = ~pi7;
  wire tmp4967;
  assign tmp4967 = (tmp4964 & tmp4965) | (tmp4964 & tmp4966) | (tmp4965 & tmp4966);
  wire tmp4968;
  assign tmp4968 = ~pi6;
  wire tmp4969;
  assign tmp4969 = 1'b1;
  wire tmp4970;
  assign tmp4970 = 1'b1;
  wire tmp4971;
  assign tmp4971 = (tmp4968 & tmp4969) | (tmp4968 & tmp4970) | (tmp4969 & tmp4970);
  wire tmp4972;
  assign tmp4972 = ~pi7;
  wire tmp4973;
  assign tmp4973 = 1'b1;
  wire tmp4974;
  assign tmp4974 = 1'b0;
  wire tmp4975;
  assign tmp4975 = (tmp4972 & tmp4973) | (tmp4972 & tmp4974) | (tmp4973 & tmp4974);
  wire tmp4976;
  assign tmp4976 = (tmp4967 & tmp4971) | (tmp4967 & tmp4975) | (tmp4971 & tmp4975);
  wire tmp4977;
  assign tmp4977 = (tmp4950 & tmp4963) | (tmp4950 & tmp4976) | (tmp4963 & tmp4976);
  wire tmp4978;
  assign tmp4978 = (tmp4897 & tmp4937) | (tmp4897 & tmp4977) | (tmp4937 & tmp4977);
  wire tmp4979;
  assign tmp4979 = 1'b0;
  wire tmp4980;
  assign tmp4980 = 1'b1;
  wire tmp4981;
  assign tmp4981 = 1'b0;
  wire tmp4982;
  assign tmp4982 = (tmp4979 & tmp4980) | (tmp4979 & tmp4981) | (tmp4980 & tmp4981);
  wire tmp4983;
  assign tmp4983 = 1'b1;
  wire tmp4984;
  assign tmp4984 = 1'b1;
  wire tmp4985;
  assign tmp4985 = 1'b1;
  wire tmp4986;
  assign tmp4986 = (tmp4983 & tmp4984) | (tmp4983 & tmp4985) | (tmp4984 & tmp4985);
  wire tmp4987;
  assign tmp4987 = 1'b0;
  wire tmp4988;
  assign tmp4988 = 1'b1;
  wire tmp4989;
  assign tmp4989 = 1'b0;
  wire tmp4990;
  assign tmp4990 = (tmp4987 & tmp4988) | (tmp4987 & tmp4989) | (tmp4988 & tmp4989);
  wire tmp4991;
  assign tmp4991 = (tmp4982 & tmp4986) | (tmp4982 & tmp4990) | (tmp4986 & tmp4990);
  wire tmp4992;
  assign tmp4992 = 1'b1;
  wire tmp4993;
  assign tmp4993 = 1'b1;
  wire tmp4994;
  assign tmp4994 = 1'b1;
  wire tmp4995;
  assign tmp4995 = (tmp4992 & tmp4993) | (tmp4992 & tmp4994) | (tmp4993 & tmp4994);
  wire tmp4996;
  assign tmp4996 = 1'b1;
  wire tmp4997;
  assign tmp4997 = ~pi5;
  wire tmp4998;
  assign tmp4998 = ~pi6;
  wire tmp4999;
  assign tmp4999 = (tmp4996 & tmp4997) | (tmp4996 & tmp4998) | (tmp4997 & tmp4998);
  wire tmp5000;
  assign tmp5000 = 1'b1;
  wire tmp5001;
  assign tmp5001 = ~pi6;
  wire tmp5002;
  assign tmp5002 = ~pi7;
  wire tmp5003;
  assign tmp5003 = (tmp5000 & tmp5001) | (tmp5000 & tmp5002) | (tmp5001 & tmp5002);
  wire tmp5004;
  assign tmp5004 = (tmp4995 & tmp4999) | (tmp4995 & tmp5003) | (tmp4999 & tmp5003);
  wire tmp5005;
  assign tmp5005 = 1'b0;
  wire tmp5006;
  assign tmp5006 = 1'b1;
  wire tmp5007;
  assign tmp5007 = 1'b0;
  wire tmp5008;
  assign tmp5008 = (tmp5005 & tmp5006) | (tmp5005 & tmp5007) | (tmp5006 & tmp5007);
  wire tmp5009;
  assign tmp5009 = 1'b1;
  wire tmp5010;
  assign tmp5010 = ~pi6;
  wire tmp5011;
  assign tmp5011 = ~pi7;
  wire tmp5012;
  assign tmp5012 = (tmp5009 & tmp5010) | (tmp5009 & tmp5011) | (tmp5010 & tmp5011);
  wire tmp5013;
  assign tmp5013 = 1'b0;
  wire tmp5014;
  assign tmp5014 = ~pi7;
  wire tmp5015;
  assign tmp5015 = 1'b0;
  wire tmp5016;
  assign tmp5016 = (tmp5013 & tmp5014) | (tmp5013 & tmp5015) | (tmp5014 & tmp5015);
  wire tmp5017;
  assign tmp5017 = (tmp5008 & tmp5012) | (tmp5008 & tmp5016) | (tmp5012 & tmp5016);
  wire tmp5018;
  assign tmp5018 = (tmp4991 & tmp5004) | (tmp4991 & tmp5017) | (tmp5004 & tmp5017);
  wire tmp5019;
  assign tmp5019 = 1'b1;
  wire tmp5020;
  assign tmp5020 = 1'b1;
  wire tmp5021;
  assign tmp5021 = 1'b1;
  wire tmp5022;
  assign tmp5022 = (tmp5019 & tmp5020) | (tmp5019 & tmp5021) | (tmp5020 & tmp5021);
  wire tmp5023;
  assign tmp5023 = 1'b1;
  wire tmp5024;
  assign tmp5024 = ~pi5;
  wire tmp5025;
  assign tmp5025 = ~pi6;
  wire tmp5026;
  assign tmp5026 = (tmp5023 & tmp5024) | (tmp5023 & tmp5025) | (tmp5024 & tmp5025);
  wire tmp5027;
  assign tmp5027 = 1'b1;
  wire tmp5028;
  assign tmp5028 = ~pi6;
  wire tmp5029;
  assign tmp5029 = ~pi7;
  wire tmp5030;
  assign tmp5030 = (tmp5027 & tmp5028) | (tmp5027 & tmp5029) | (tmp5028 & tmp5029);
  wire tmp5031;
  assign tmp5031 = (tmp5022 & tmp5026) | (tmp5022 & tmp5030) | (tmp5026 & tmp5030);
  wire tmp5032;
  assign tmp5032 = 1'b1;
  wire tmp5033;
  assign tmp5033 = ~pi5;
  wire tmp5034;
  assign tmp5034 = ~pi6;
  wire tmp5035;
  assign tmp5035 = (tmp5032 & tmp5033) | (tmp5032 & tmp5034) | (tmp5033 & tmp5034);
  wire tmp5036;
  assign tmp5036 = ~pi5;
  wire tmp5037;
  assign tmp5037 = 1'b1;
  wire tmp5038;
  assign tmp5038 = 1'b1;
  wire tmp5039;
  assign tmp5039 = (tmp5036 & tmp5037) | (tmp5036 & tmp5038) | (tmp5037 & tmp5038);
  wire tmp5040;
  assign tmp5040 = ~pi6;
  wire tmp5041;
  assign tmp5041 = 1'b1;
  wire tmp5042;
  assign tmp5042 = 1'b1;
  wire tmp5043;
  assign tmp5043 = (tmp5040 & tmp5041) | (tmp5040 & tmp5042) | (tmp5041 & tmp5042);
  wire tmp5044;
  assign tmp5044 = (tmp5035 & tmp5039) | (tmp5035 & tmp5043) | (tmp5039 & tmp5043);
  wire tmp5045;
  assign tmp5045 = 1'b1;
  wire tmp5046;
  assign tmp5046 = ~pi6;
  wire tmp5047;
  assign tmp5047 = ~pi7;
  wire tmp5048;
  assign tmp5048 = (tmp5045 & tmp5046) | (tmp5045 & tmp5047) | (tmp5046 & tmp5047);
  wire tmp5049;
  assign tmp5049 = ~pi6;
  wire tmp5050;
  assign tmp5050 = 1'b1;
  wire tmp5051;
  assign tmp5051 = 1'b1;
  wire tmp5052;
  assign tmp5052 = (tmp5049 & tmp5050) | (tmp5049 & tmp5051) | (tmp5050 & tmp5051);
  wire tmp5053;
  assign tmp5053 = ~pi7;
  wire tmp5054;
  assign tmp5054 = 1'b1;
  wire tmp5055;
  assign tmp5055 = 1'b0;
  wire tmp5056;
  assign tmp5056 = (tmp5053 & tmp5054) | (tmp5053 & tmp5055) | (tmp5054 & tmp5055);
  wire tmp5057;
  assign tmp5057 = (tmp5048 & tmp5052) | (tmp5048 & tmp5056) | (tmp5052 & tmp5056);
  wire tmp5058;
  assign tmp5058 = (tmp5031 & tmp5044) | (tmp5031 & tmp5057) | (tmp5044 & tmp5057);
  wire tmp5059;
  assign tmp5059 = 1'b0;
  wire tmp5060;
  assign tmp5060 = 1'b1;
  wire tmp5061;
  assign tmp5061 = 1'b0;
  wire tmp5062;
  assign tmp5062 = (tmp5059 & tmp5060) | (tmp5059 & tmp5061) | (tmp5060 & tmp5061);
  wire tmp5063;
  assign tmp5063 = 1'b1;
  wire tmp5064;
  assign tmp5064 = ~pi6;
  wire tmp5065;
  assign tmp5065 = ~pi7;
  wire tmp5066;
  assign tmp5066 = (tmp5063 & tmp5064) | (tmp5063 & tmp5065) | (tmp5064 & tmp5065);
  wire tmp5067;
  assign tmp5067 = 1'b0;
  wire tmp5068;
  assign tmp5068 = ~pi7;
  wire tmp5069;
  assign tmp5069 = 1'b0;
  wire tmp5070;
  assign tmp5070 = (tmp5067 & tmp5068) | (tmp5067 & tmp5069) | (tmp5068 & tmp5069);
  wire tmp5071;
  assign tmp5071 = (tmp5062 & tmp5066) | (tmp5062 & tmp5070) | (tmp5066 & tmp5070);
  wire tmp5072;
  assign tmp5072 = 1'b1;
  wire tmp5073;
  assign tmp5073 = ~pi6;
  wire tmp5074;
  assign tmp5074 = ~pi7;
  wire tmp5075;
  assign tmp5075 = (tmp5072 & tmp5073) | (tmp5072 & tmp5074) | (tmp5073 & tmp5074);
  wire tmp5076;
  assign tmp5076 = ~pi6;
  wire tmp5077;
  assign tmp5077 = 1'b1;
  wire tmp5078;
  assign tmp5078 = 1'b1;
  wire tmp5079;
  assign tmp5079 = (tmp5076 & tmp5077) | (tmp5076 & tmp5078) | (tmp5077 & tmp5078);
  wire tmp5080;
  assign tmp5080 = ~pi7;
  wire tmp5081;
  assign tmp5081 = 1'b1;
  wire tmp5082;
  assign tmp5082 = 1'b0;
  wire tmp5083;
  assign tmp5083 = (tmp5080 & tmp5081) | (tmp5080 & tmp5082) | (tmp5081 & tmp5082);
  wire tmp5084;
  assign tmp5084 = (tmp5075 & tmp5079) | (tmp5075 & tmp5083) | (tmp5079 & tmp5083);
  wire tmp5085;
  assign tmp5085 = 1'b0;
  wire tmp5086;
  assign tmp5086 = ~pi7;
  wire tmp5087;
  assign tmp5087 = 1'b0;
  wire tmp5088;
  assign tmp5088 = (tmp5085 & tmp5086) | (tmp5085 & tmp5087) | (tmp5086 & tmp5087);
  wire tmp5089;
  assign tmp5089 = ~pi7;
  wire tmp5090;
  assign tmp5090 = 1'b1;
  wire tmp5091;
  assign tmp5091 = 1'b0;
  wire tmp5092;
  assign tmp5092 = (tmp5089 & tmp5090) | (tmp5089 & tmp5091) | (tmp5090 & tmp5091);
  wire tmp5093;
  assign tmp5093 = 1'b0;
  wire tmp5094;
  assign tmp5094 = 1'b0;
  wire tmp5095;
  assign tmp5095 = 1'b0;
  wire tmp5096;
  assign tmp5096 = (tmp5093 & tmp5094) | (tmp5093 & tmp5095) | (tmp5094 & tmp5095);
  wire tmp5097;
  assign tmp5097 = (tmp5088 & tmp5092) | (tmp5088 & tmp5096) | (tmp5092 & tmp5096);
  wire tmp5098;
  assign tmp5098 = (tmp5071 & tmp5084) | (tmp5071 & tmp5097) | (tmp5084 & tmp5097);
  wire tmp5099;
  assign tmp5099 = (tmp5018 & tmp5058) | (tmp5018 & tmp5098) | (tmp5058 & tmp5098);
  wire tmp5100;
  assign tmp5100 = (tmp4857 & tmp4978) | (tmp4857 & tmp5099) | (tmp4978 & tmp5099);
  wire tmp5101;
  assign tmp5101 = 1'b0;
  wire tmp5102;
  assign tmp5102 = 1'b0;
  wire tmp5103;
  assign tmp5103 = 1'b0;
  wire tmp5104;
  assign tmp5104 = (tmp5101 & tmp5102) | (tmp5101 & tmp5103) | (tmp5102 & tmp5103);
  wire tmp5105;
  assign tmp5105 = 1'b0;
  wire tmp5106;
  assign tmp5106 = 1'b1;
  wire tmp5107;
  assign tmp5107 = 1'b0;
  wire tmp5108;
  assign tmp5108 = (tmp5105 & tmp5106) | (tmp5105 & tmp5107) | (tmp5106 & tmp5107);
  wire tmp5109;
  assign tmp5109 = 1'b0;
  wire tmp5110;
  assign tmp5110 = 1'b0;
  wire tmp5111;
  assign tmp5111 = 1'b0;
  wire tmp5112;
  assign tmp5112 = (tmp5109 & tmp5110) | (tmp5109 & tmp5111) | (tmp5110 & tmp5111);
  wire tmp5113;
  assign tmp5113 = (tmp5104 & tmp5108) | (tmp5104 & tmp5112) | (tmp5108 & tmp5112);
  wire tmp5114;
  assign tmp5114 = 1'b0;
  wire tmp5115;
  assign tmp5115 = 1'b1;
  wire tmp5116;
  assign tmp5116 = 1'b0;
  wire tmp5117;
  assign tmp5117 = (tmp5114 & tmp5115) | (tmp5114 & tmp5116) | (tmp5115 & tmp5116);
  wire tmp5118;
  assign tmp5118 = 1'b1;
  wire tmp5119;
  assign tmp5119 = 1'b1;
  wire tmp5120;
  assign tmp5120 = 1'b1;
  wire tmp5121;
  assign tmp5121 = (tmp5118 & tmp5119) | (tmp5118 & tmp5120) | (tmp5119 & tmp5120);
  wire tmp5122;
  assign tmp5122 = 1'b0;
  wire tmp5123;
  assign tmp5123 = 1'b1;
  wire tmp5124;
  assign tmp5124 = 1'b0;
  wire tmp5125;
  assign tmp5125 = (tmp5122 & tmp5123) | (tmp5122 & tmp5124) | (tmp5123 & tmp5124);
  wire tmp5126;
  assign tmp5126 = (tmp5117 & tmp5121) | (tmp5117 & tmp5125) | (tmp5121 & tmp5125);
  wire tmp5127;
  assign tmp5127 = 1'b0;
  wire tmp5128;
  assign tmp5128 = 1'b0;
  wire tmp5129;
  assign tmp5129 = 1'b0;
  wire tmp5130;
  assign tmp5130 = (tmp5127 & tmp5128) | (tmp5127 & tmp5129) | (tmp5128 & tmp5129);
  wire tmp5131;
  assign tmp5131 = 1'b0;
  wire tmp5132;
  assign tmp5132 = 1'b1;
  wire tmp5133;
  assign tmp5133 = 1'b0;
  wire tmp5134;
  assign tmp5134 = (tmp5131 & tmp5132) | (tmp5131 & tmp5133) | (tmp5132 & tmp5133);
  wire tmp5135;
  assign tmp5135 = 1'b0;
  wire tmp5136;
  assign tmp5136 = 1'b0;
  wire tmp5137;
  assign tmp5137 = 1'b0;
  wire tmp5138;
  assign tmp5138 = (tmp5135 & tmp5136) | (tmp5135 & tmp5137) | (tmp5136 & tmp5137);
  wire tmp5139;
  assign tmp5139 = (tmp5130 & tmp5134) | (tmp5130 & tmp5138) | (tmp5134 & tmp5138);
  wire tmp5140;
  assign tmp5140 = (tmp5113 & tmp5126) | (tmp5113 & tmp5139) | (tmp5126 & tmp5139);
  wire tmp5141;
  assign tmp5141 = 1'b0;
  wire tmp5142;
  assign tmp5142 = 1'b1;
  wire tmp5143;
  assign tmp5143 = 1'b0;
  wire tmp5144;
  assign tmp5144 = (tmp5141 & tmp5142) | (tmp5141 & tmp5143) | (tmp5142 & tmp5143);
  wire tmp5145;
  assign tmp5145 = 1'b1;
  wire tmp5146;
  assign tmp5146 = 1'b1;
  wire tmp5147;
  assign tmp5147 = 1'b1;
  wire tmp5148;
  assign tmp5148 = (tmp5145 & tmp5146) | (tmp5145 & tmp5147) | (tmp5146 & tmp5147);
  wire tmp5149;
  assign tmp5149 = 1'b0;
  wire tmp5150;
  assign tmp5150 = 1'b1;
  wire tmp5151;
  assign tmp5151 = 1'b0;
  wire tmp5152;
  assign tmp5152 = (tmp5149 & tmp5150) | (tmp5149 & tmp5151) | (tmp5150 & tmp5151);
  wire tmp5153;
  assign tmp5153 = (tmp5144 & tmp5148) | (tmp5144 & tmp5152) | (tmp5148 & tmp5152);
  wire tmp5154;
  assign tmp5154 = 1'b1;
  wire tmp5155;
  assign tmp5155 = 1'b1;
  wire tmp5156;
  assign tmp5156 = 1'b1;
  wire tmp5157;
  assign tmp5157 = (tmp5154 & tmp5155) | (tmp5154 & tmp5156) | (tmp5155 & tmp5156);
  wire tmp5158;
  assign tmp5158 = 1'b1;
  wire tmp5159;
  assign tmp5159 = ~pi5;
  wire tmp5160;
  assign tmp5160 = ~pi6;
  wire tmp5161;
  assign tmp5161 = (tmp5158 & tmp5159) | (tmp5158 & tmp5160) | (tmp5159 & tmp5160);
  wire tmp5162;
  assign tmp5162 = 1'b1;
  wire tmp5163;
  assign tmp5163 = ~pi6;
  wire tmp5164;
  assign tmp5164 = ~pi7;
  wire tmp5165;
  assign tmp5165 = (tmp5162 & tmp5163) | (tmp5162 & tmp5164) | (tmp5163 & tmp5164);
  wire tmp5166;
  assign tmp5166 = (tmp5157 & tmp5161) | (tmp5157 & tmp5165) | (tmp5161 & tmp5165);
  wire tmp5167;
  assign tmp5167 = 1'b0;
  wire tmp5168;
  assign tmp5168 = 1'b1;
  wire tmp5169;
  assign tmp5169 = 1'b0;
  wire tmp5170;
  assign tmp5170 = (tmp5167 & tmp5168) | (tmp5167 & tmp5169) | (tmp5168 & tmp5169);
  wire tmp5171;
  assign tmp5171 = 1'b1;
  wire tmp5172;
  assign tmp5172 = ~pi6;
  wire tmp5173;
  assign tmp5173 = ~pi7;
  wire tmp5174;
  assign tmp5174 = (tmp5171 & tmp5172) | (tmp5171 & tmp5173) | (tmp5172 & tmp5173);
  wire tmp5175;
  assign tmp5175 = 1'b0;
  wire tmp5176;
  assign tmp5176 = ~pi7;
  wire tmp5177;
  assign tmp5177 = 1'b0;
  wire tmp5178;
  assign tmp5178 = (tmp5175 & tmp5176) | (tmp5175 & tmp5177) | (tmp5176 & tmp5177);
  wire tmp5179;
  assign tmp5179 = (tmp5170 & tmp5174) | (tmp5170 & tmp5178) | (tmp5174 & tmp5178);
  wire tmp5180;
  assign tmp5180 = (tmp5153 & tmp5166) | (tmp5153 & tmp5179) | (tmp5166 & tmp5179);
  wire tmp5181;
  assign tmp5181 = 1'b0;
  wire tmp5182;
  assign tmp5182 = 1'b0;
  wire tmp5183;
  assign tmp5183 = 1'b0;
  wire tmp5184;
  assign tmp5184 = (tmp5181 & tmp5182) | (tmp5181 & tmp5183) | (tmp5182 & tmp5183);
  wire tmp5185;
  assign tmp5185 = 1'b0;
  wire tmp5186;
  assign tmp5186 = 1'b1;
  wire tmp5187;
  assign tmp5187 = 1'b0;
  wire tmp5188;
  assign tmp5188 = (tmp5185 & tmp5186) | (tmp5185 & tmp5187) | (tmp5186 & tmp5187);
  wire tmp5189;
  assign tmp5189 = 1'b0;
  wire tmp5190;
  assign tmp5190 = 1'b0;
  wire tmp5191;
  assign tmp5191 = 1'b0;
  wire tmp5192;
  assign tmp5192 = (tmp5189 & tmp5190) | (tmp5189 & tmp5191) | (tmp5190 & tmp5191);
  wire tmp5193;
  assign tmp5193 = (tmp5184 & tmp5188) | (tmp5184 & tmp5192) | (tmp5188 & tmp5192);
  wire tmp5194;
  assign tmp5194 = 1'b0;
  wire tmp5195;
  assign tmp5195 = 1'b1;
  wire tmp5196;
  assign tmp5196 = 1'b0;
  wire tmp5197;
  assign tmp5197 = (tmp5194 & tmp5195) | (tmp5194 & tmp5196) | (tmp5195 & tmp5196);
  wire tmp5198;
  assign tmp5198 = 1'b1;
  wire tmp5199;
  assign tmp5199 = ~pi6;
  wire tmp5200;
  assign tmp5200 = ~pi7;
  wire tmp5201;
  assign tmp5201 = (tmp5198 & tmp5199) | (tmp5198 & tmp5200) | (tmp5199 & tmp5200);
  wire tmp5202;
  assign tmp5202 = 1'b0;
  wire tmp5203;
  assign tmp5203 = ~pi7;
  wire tmp5204;
  assign tmp5204 = 1'b0;
  wire tmp5205;
  assign tmp5205 = (tmp5202 & tmp5203) | (tmp5202 & tmp5204) | (tmp5203 & tmp5204);
  wire tmp5206;
  assign tmp5206 = (tmp5197 & tmp5201) | (tmp5197 & tmp5205) | (tmp5201 & tmp5205);
  wire tmp5207;
  assign tmp5207 = 1'b0;
  wire tmp5208;
  assign tmp5208 = 1'b0;
  wire tmp5209;
  assign tmp5209 = 1'b0;
  wire tmp5210;
  assign tmp5210 = (tmp5207 & tmp5208) | (tmp5207 & tmp5209) | (tmp5208 & tmp5209);
  wire tmp5211;
  assign tmp5211 = 1'b0;
  wire tmp5212;
  assign tmp5212 = ~pi7;
  wire tmp5213;
  assign tmp5213 = 1'b0;
  wire tmp5214;
  assign tmp5214 = (tmp5211 & tmp5212) | (tmp5211 & tmp5213) | (tmp5212 & tmp5213);
  wire tmp5215;
  assign tmp5215 = 1'b0;
  wire tmp5216;
  assign tmp5216 = 1'b0;
  wire tmp5217;
  assign tmp5217 = 1'b0;
  wire tmp5218;
  assign tmp5218 = (tmp5215 & tmp5216) | (tmp5215 & tmp5217) | (tmp5216 & tmp5217);
  wire tmp5219;
  assign tmp5219 = (tmp5210 & tmp5214) | (tmp5210 & tmp5218) | (tmp5214 & tmp5218);
  wire tmp5220;
  assign tmp5220 = (tmp5193 & tmp5206) | (tmp5193 & tmp5219) | (tmp5206 & tmp5219);
  wire tmp5221;
  assign tmp5221 = (tmp5140 & tmp5180) | (tmp5140 & tmp5220) | (tmp5180 & tmp5220);
  wire tmp5222;
  assign tmp5222 = 1'b0;
  wire tmp5223;
  assign tmp5223 = 1'b1;
  wire tmp5224;
  assign tmp5224 = 1'b0;
  wire tmp5225;
  assign tmp5225 = (tmp5222 & tmp5223) | (tmp5222 & tmp5224) | (tmp5223 & tmp5224);
  wire tmp5226;
  assign tmp5226 = 1'b1;
  wire tmp5227;
  assign tmp5227 = 1'b1;
  wire tmp5228;
  assign tmp5228 = 1'b1;
  wire tmp5229;
  assign tmp5229 = (tmp5226 & tmp5227) | (tmp5226 & tmp5228) | (tmp5227 & tmp5228);
  wire tmp5230;
  assign tmp5230 = 1'b0;
  wire tmp5231;
  assign tmp5231 = 1'b1;
  wire tmp5232;
  assign tmp5232 = 1'b0;
  wire tmp5233;
  assign tmp5233 = (tmp5230 & tmp5231) | (tmp5230 & tmp5232) | (tmp5231 & tmp5232);
  wire tmp5234;
  assign tmp5234 = (tmp5225 & tmp5229) | (tmp5225 & tmp5233) | (tmp5229 & tmp5233);
  wire tmp5235;
  assign tmp5235 = 1'b1;
  wire tmp5236;
  assign tmp5236 = 1'b1;
  wire tmp5237;
  assign tmp5237 = 1'b1;
  wire tmp5238;
  assign tmp5238 = (tmp5235 & tmp5236) | (tmp5235 & tmp5237) | (tmp5236 & tmp5237);
  wire tmp5239;
  assign tmp5239 = 1'b1;
  wire tmp5240;
  assign tmp5240 = ~pi5;
  wire tmp5241;
  assign tmp5241 = ~pi6;
  wire tmp5242;
  assign tmp5242 = (tmp5239 & tmp5240) | (tmp5239 & tmp5241) | (tmp5240 & tmp5241);
  wire tmp5243;
  assign tmp5243 = 1'b1;
  wire tmp5244;
  assign tmp5244 = ~pi6;
  wire tmp5245;
  assign tmp5245 = ~pi7;
  wire tmp5246;
  assign tmp5246 = (tmp5243 & tmp5244) | (tmp5243 & tmp5245) | (tmp5244 & tmp5245);
  wire tmp5247;
  assign tmp5247 = (tmp5238 & tmp5242) | (tmp5238 & tmp5246) | (tmp5242 & tmp5246);
  wire tmp5248;
  assign tmp5248 = 1'b0;
  wire tmp5249;
  assign tmp5249 = 1'b1;
  wire tmp5250;
  assign tmp5250 = 1'b0;
  wire tmp5251;
  assign tmp5251 = (tmp5248 & tmp5249) | (tmp5248 & tmp5250) | (tmp5249 & tmp5250);
  wire tmp5252;
  assign tmp5252 = 1'b1;
  wire tmp5253;
  assign tmp5253 = ~pi6;
  wire tmp5254;
  assign tmp5254 = ~pi7;
  wire tmp5255;
  assign tmp5255 = (tmp5252 & tmp5253) | (tmp5252 & tmp5254) | (tmp5253 & tmp5254);
  wire tmp5256;
  assign tmp5256 = 1'b0;
  wire tmp5257;
  assign tmp5257 = ~pi7;
  wire tmp5258;
  assign tmp5258 = 1'b0;
  wire tmp5259;
  assign tmp5259 = (tmp5256 & tmp5257) | (tmp5256 & tmp5258) | (tmp5257 & tmp5258);
  wire tmp5260;
  assign tmp5260 = (tmp5251 & tmp5255) | (tmp5251 & tmp5259) | (tmp5255 & tmp5259);
  wire tmp5261;
  assign tmp5261 = (tmp5234 & tmp5247) | (tmp5234 & tmp5260) | (tmp5247 & tmp5260);
  wire tmp5262;
  assign tmp5262 = 1'b1;
  wire tmp5263;
  assign tmp5263 = 1'b1;
  wire tmp5264;
  assign tmp5264 = 1'b1;
  wire tmp5265;
  assign tmp5265 = (tmp5262 & tmp5263) | (tmp5262 & tmp5264) | (tmp5263 & tmp5264);
  wire tmp5266;
  assign tmp5266 = 1'b1;
  wire tmp5267;
  assign tmp5267 = ~pi5;
  wire tmp5268;
  assign tmp5268 = ~pi6;
  wire tmp5269;
  assign tmp5269 = (tmp5266 & tmp5267) | (tmp5266 & tmp5268) | (tmp5267 & tmp5268);
  wire tmp5270;
  assign tmp5270 = 1'b1;
  wire tmp5271;
  assign tmp5271 = ~pi6;
  wire tmp5272;
  assign tmp5272 = ~pi7;
  wire tmp5273;
  assign tmp5273 = (tmp5270 & tmp5271) | (tmp5270 & tmp5272) | (tmp5271 & tmp5272);
  wire tmp5274;
  assign tmp5274 = (tmp5265 & tmp5269) | (tmp5265 & tmp5273) | (tmp5269 & tmp5273);
  wire tmp5275;
  assign tmp5275 = 1'b1;
  wire tmp5276;
  assign tmp5276 = ~pi5;
  wire tmp5277;
  assign tmp5277 = ~pi6;
  wire tmp5278;
  assign tmp5278 = (tmp5275 & tmp5276) | (tmp5275 & tmp5277) | (tmp5276 & tmp5277);
  wire tmp5279;
  assign tmp5279 = ~pi5;
  wire tmp5280;
  assign tmp5280 = 1'b1;
  wire tmp5281;
  assign tmp5281 = 1'b1;
  wire tmp5282;
  assign tmp5282 = (tmp5279 & tmp5280) | (tmp5279 & tmp5281) | (tmp5280 & tmp5281);
  wire tmp5283;
  assign tmp5283 = ~pi6;
  wire tmp5284;
  assign tmp5284 = 1'b1;
  wire tmp5285;
  assign tmp5285 = 1'b1;
  wire tmp5286;
  assign tmp5286 = (tmp5283 & tmp5284) | (tmp5283 & tmp5285) | (tmp5284 & tmp5285);
  wire tmp5287;
  assign tmp5287 = (tmp5278 & tmp5282) | (tmp5278 & tmp5286) | (tmp5282 & tmp5286);
  wire tmp5288;
  assign tmp5288 = 1'b1;
  wire tmp5289;
  assign tmp5289 = ~pi6;
  wire tmp5290;
  assign tmp5290 = ~pi7;
  wire tmp5291;
  assign tmp5291 = (tmp5288 & tmp5289) | (tmp5288 & tmp5290) | (tmp5289 & tmp5290);
  wire tmp5292;
  assign tmp5292 = ~pi6;
  wire tmp5293;
  assign tmp5293 = 1'b1;
  wire tmp5294;
  assign tmp5294 = 1'b1;
  wire tmp5295;
  assign tmp5295 = (tmp5292 & tmp5293) | (tmp5292 & tmp5294) | (tmp5293 & tmp5294);
  wire tmp5296;
  assign tmp5296 = ~pi7;
  wire tmp5297;
  assign tmp5297 = 1'b1;
  wire tmp5298;
  assign tmp5298 = 1'b0;
  wire tmp5299;
  assign tmp5299 = (tmp5296 & tmp5297) | (tmp5296 & tmp5298) | (tmp5297 & tmp5298);
  wire tmp5300;
  assign tmp5300 = (tmp5291 & tmp5295) | (tmp5291 & tmp5299) | (tmp5295 & tmp5299);
  wire tmp5301;
  assign tmp5301 = (tmp5274 & tmp5287) | (tmp5274 & tmp5300) | (tmp5287 & tmp5300);
  wire tmp5302;
  assign tmp5302 = 1'b0;
  wire tmp5303;
  assign tmp5303 = 1'b1;
  wire tmp5304;
  assign tmp5304 = 1'b0;
  wire tmp5305;
  assign tmp5305 = (tmp5302 & tmp5303) | (tmp5302 & tmp5304) | (tmp5303 & tmp5304);
  wire tmp5306;
  assign tmp5306 = 1'b1;
  wire tmp5307;
  assign tmp5307 = ~pi6;
  wire tmp5308;
  assign tmp5308 = ~pi7;
  wire tmp5309;
  assign tmp5309 = (tmp5306 & tmp5307) | (tmp5306 & tmp5308) | (tmp5307 & tmp5308);
  wire tmp5310;
  assign tmp5310 = 1'b0;
  wire tmp5311;
  assign tmp5311 = ~pi7;
  wire tmp5312;
  assign tmp5312 = 1'b0;
  wire tmp5313;
  assign tmp5313 = (tmp5310 & tmp5311) | (tmp5310 & tmp5312) | (tmp5311 & tmp5312);
  wire tmp5314;
  assign tmp5314 = (tmp5305 & tmp5309) | (tmp5305 & tmp5313) | (tmp5309 & tmp5313);
  wire tmp5315;
  assign tmp5315 = 1'b1;
  wire tmp5316;
  assign tmp5316 = ~pi6;
  wire tmp5317;
  assign tmp5317 = ~pi7;
  wire tmp5318;
  assign tmp5318 = (tmp5315 & tmp5316) | (tmp5315 & tmp5317) | (tmp5316 & tmp5317);
  wire tmp5319;
  assign tmp5319 = ~pi6;
  wire tmp5320;
  assign tmp5320 = 1'b1;
  wire tmp5321;
  assign tmp5321 = 1'b1;
  wire tmp5322;
  assign tmp5322 = (tmp5319 & tmp5320) | (tmp5319 & tmp5321) | (tmp5320 & tmp5321);
  wire tmp5323;
  assign tmp5323 = ~pi7;
  wire tmp5324;
  assign tmp5324 = 1'b1;
  wire tmp5325;
  assign tmp5325 = 1'b0;
  wire tmp5326;
  assign tmp5326 = (tmp5323 & tmp5324) | (tmp5323 & tmp5325) | (tmp5324 & tmp5325);
  wire tmp5327;
  assign tmp5327 = (tmp5318 & tmp5322) | (tmp5318 & tmp5326) | (tmp5322 & tmp5326);
  wire tmp5328;
  assign tmp5328 = 1'b0;
  wire tmp5329;
  assign tmp5329 = ~pi7;
  wire tmp5330;
  assign tmp5330 = 1'b0;
  wire tmp5331;
  assign tmp5331 = (tmp5328 & tmp5329) | (tmp5328 & tmp5330) | (tmp5329 & tmp5330);
  wire tmp5332;
  assign tmp5332 = ~pi7;
  wire tmp5333;
  assign tmp5333 = 1'b1;
  wire tmp5334;
  assign tmp5334 = 1'b0;
  wire tmp5335;
  assign tmp5335 = (tmp5332 & tmp5333) | (tmp5332 & tmp5334) | (tmp5333 & tmp5334);
  wire tmp5336;
  assign tmp5336 = 1'b0;
  wire tmp5337;
  assign tmp5337 = 1'b0;
  wire tmp5338;
  assign tmp5338 = 1'b0;
  wire tmp5339;
  assign tmp5339 = (tmp5336 & tmp5337) | (tmp5336 & tmp5338) | (tmp5337 & tmp5338);
  wire tmp5340;
  assign tmp5340 = (tmp5331 & tmp5335) | (tmp5331 & tmp5339) | (tmp5335 & tmp5339);
  wire tmp5341;
  assign tmp5341 = (tmp5314 & tmp5327) | (tmp5314 & tmp5340) | (tmp5327 & tmp5340);
  wire tmp5342;
  assign tmp5342 = (tmp5261 & tmp5301) | (tmp5261 & tmp5341) | (tmp5301 & tmp5341);
  wire tmp5343;
  assign tmp5343 = 1'b0;
  wire tmp5344;
  assign tmp5344 = 1'b0;
  wire tmp5345;
  assign tmp5345 = 1'b0;
  wire tmp5346;
  assign tmp5346 = (tmp5343 & tmp5344) | (tmp5343 & tmp5345) | (tmp5344 & tmp5345);
  wire tmp5347;
  assign tmp5347 = 1'b0;
  wire tmp5348;
  assign tmp5348 = 1'b1;
  wire tmp5349;
  assign tmp5349 = 1'b0;
  wire tmp5350;
  assign tmp5350 = (tmp5347 & tmp5348) | (tmp5347 & tmp5349) | (tmp5348 & tmp5349);
  wire tmp5351;
  assign tmp5351 = 1'b0;
  wire tmp5352;
  assign tmp5352 = 1'b0;
  wire tmp5353;
  assign tmp5353 = 1'b0;
  wire tmp5354;
  assign tmp5354 = (tmp5351 & tmp5352) | (tmp5351 & tmp5353) | (tmp5352 & tmp5353);
  wire tmp5355;
  assign tmp5355 = (tmp5346 & tmp5350) | (tmp5346 & tmp5354) | (tmp5350 & tmp5354);
  wire tmp5356;
  assign tmp5356 = 1'b0;
  wire tmp5357;
  assign tmp5357 = 1'b1;
  wire tmp5358;
  assign tmp5358 = 1'b0;
  wire tmp5359;
  assign tmp5359 = (tmp5356 & tmp5357) | (tmp5356 & tmp5358) | (tmp5357 & tmp5358);
  wire tmp5360;
  assign tmp5360 = 1'b1;
  wire tmp5361;
  assign tmp5361 = ~pi6;
  wire tmp5362;
  assign tmp5362 = ~pi7;
  wire tmp5363;
  assign tmp5363 = (tmp5360 & tmp5361) | (tmp5360 & tmp5362) | (tmp5361 & tmp5362);
  wire tmp5364;
  assign tmp5364 = 1'b0;
  wire tmp5365;
  assign tmp5365 = ~pi7;
  wire tmp5366;
  assign tmp5366 = 1'b0;
  wire tmp5367;
  assign tmp5367 = (tmp5364 & tmp5365) | (tmp5364 & tmp5366) | (tmp5365 & tmp5366);
  wire tmp5368;
  assign tmp5368 = (tmp5359 & tmp5363) | (tmp5359 & tmp5367) | (tmp5363 & tmp5367);
  wire tmp5369;
  assign tmp5369 = 1'b0;
  wire tmp5370;
  assign tmp5370 = 1'b0;
  wire tmp5371;
  assign tmp5371 = 1'b0;
  wire tmp5372;
  assign tmp5372 = (tmp5369 & tmp5370) | (tmp5369 & tmp5371) | (tmp5370 & tmp5371);
  wire tmp5373;
  assign tmp5373 = 1'b0;
  wire tmp5374;
  assign tmp5374 = ~pi7;
  wire tmp5375;
  assign tmp5375 = 1'b0;
  wire tmp5376;
  assign tmp5376 = (tmp5373 & tmp5374) | (tmp5373 & tmp5375) | (tmp5374 & tmp5375);
  wire tmp5377;
  assign tmp5377 = 1'b0;
  wire tmp5378;
  assign tmp5378 = 1'b0;
  wire tmp5379;
  assign tmp5379 = 1'b0;
  wire tmp5380;
  assign tmp5380 = (tmp5377 & tmp5378) | (tmp5377 & tmp5379) | (tmp5378 & tmp5379);
  wire tmp5381;
  assign tmp5381 = (tmp5372 & tmp5376) | (tmp5372 & tmp5380) | (tmp5376 & tmp5380);
  wire tmp5382;
  assign tmp5382 = (tmp5355 & tmp5368) | (tmp5355 & tmp5381) | (tmp5368 & tmp5381);
  wire tmp5383;
  assign tmp5383 = 1'b0;
  wire tmp5384;
  assign tmp5384 = 1'b1;
  wire tmp5385;
  assign tmp5385 = 1'b0;
  wire tmp5386;
  assign tmp5386 = (tmp5383 & tmp5384) | (tmp5383 & tmp5385) | (tmp5384 & tmp5385);
  wire tmp5387;
  assign tmp5387 = 1'b1;
  wire tmp5388;
  assign tmp5388 = ~pi6;
  wire tmp5389;
  assign tmp5389 = ~pi7;
  wire tmp5390;
  assign tmp5390 = (tmp5387 & tmp5388) | (tmp5387 & tmp5389) | (tmp5388 & tmp5389);
  wire tmp5391;
  assign tmp5391 = 1'b0;
  wire tmp5392;
  assign tmp5392 = ~pi7;
  wire tmp5393;
  assign tmp5393 = 1'b0;
  wire tmp5394;
  assign tmp5394 = (tmp5391 & tmp5392) | (tmp5391 & tmp5393) | (tmp5392 & tmp5393);
  wire tmp5395;
  assign tmp5395 = (tmp5386 & tmp5390) | (tmp5386 & tmp5394) | (tmp5390 & tmp5394);
  wire tmp5396;
  assign tmp5396 = 1'b1;
  wire tmp5397;
  assign tmp5397 = ~pi6;
  wire tmp5398;
  assign tmp5398 = ~pi7;
  wire tmp5399;
  assign tmp5399 = (tmp5396 & tmp5397) | (tmp5396 & tmp5398) | (tmp5397 & tmp5398);
  wire tmp5400;
  assign tmp5400 = ~pi6;
  wire tmp5401;
  assign tmp5401 = 1'b1;
  wire tmp5402;
  assign tmp5402 = 1'b1;
  wire tmp5403;
  assign tmp5403 = (tmp5400 & tmp5401) | (tmp5400 & tmp5402) | (tmp5401 & tmp5402);
  wire tmp5404;
  assign tmp5404 = ~pi7;
  wire tmp5405;
  assign tmp5405 = 1'b1;
  wire tmp5406;
  assign tmp5406 = 1'b0;
  wire tmp5407;
  assign tmp5407 = (tmp5404 & tmp5405) | (tmp5404 & tmp5406) | (tmp5405 & tmp5406);
  wire tmp5408;
  assign tmp5408 = (tmp5399 & tmp5403) | (tmp5399 & tmp5407) | (tmp5403 & tmp5407);
  wire tmp5409;
  assign tmp5409 = 1'b0;
  wire tmp5410;
  assign tmp5410 = ~pi7;
  wire tmp5411;
  assign tmp5411 = 1'b0;
  wire tmp5412;
  assign tmp5412 = (tmp5409 & tmp5410) | (tmp5409 & tmp5411) | (tmp5410 & tmp5411);
  wire tmp5413;
  assign tmp5413 = ~pi7;
  wire tmp5414;
  assign tmp5414 = 1'b1;
  wire tmp5415;
  assign tmp5415 = 1'b0;
  wire tmp5416;
  assign tmp5416 = (tmp5413 & tmp5414) | (tmp5413 & tmp5415) | (tmp5414 & tmp5415);
  wire tmp5417;
  assign tmp5417 = 1'b0;
  wire tmp5418;
  assign tmp5418 = 1'b0;
  wire tmp5419;
  assign tmp5419 = 1'b0;
  wire tmp5420;
  assign tmp5420 = (tmp5417 & tmp5418) | (tmp5417 & tmp5419) | (tmp5418 & tmp5419);
  wire tmp5421;
  assign tmp5421 = (tmp5412 & tmp5416) | (tmp5412 & tmp5420) | (tmp5416 & tmp5420);
  wire tmp5422;
  assign tmp5422 = (tmp5395 & tmp5408) | (tmp5395 & tmp5421) | (tmp5408 & tmp5421);
  wire tmp5423;
  assign tmp5423 = 1'b0;
  wire tmp5424;
  assign tmp5424 = 1'b0;
  wire tmp5425;
  assign tmp5425 = 1'b0;
  wire tmp5426;
  assign tmp5426 = (tmp5423 & tmp5424) | (tmp5423 & tmp5425) | (tmp5424 & tmp5425);
  wire tmp5427;
  assign tmp5427 = 1'b0;
  wire tmp5428;
  assign tmp5428 = ~pi7;
  wire tmp5429;
  assign tmp5429 = 1'b0;
  wire tmp5430;
  assign tmp5430 = (tmp5427 & tmp5428) | (tmp5427 & tmp5429) | (tmp5428 & tmp5429);
  wire tmp5431;
  assign tmp5431 = 1'b0;
  wire tmp5432;
  assign tmp5432 = 1'b0;
  wire tmp5433;
  assign tmp5433 = 1'b0;
  wire tmp5434;
  assign tmp5434 = (tmp5431 & tmp5432) | (tmp5431 & tmp5433) | (tmp5432 & tmp5433);
  wire tmp5435;
  assign tmp5435 = (tmp5426 & tmp5430) | (tmp5426 & tmp5434) | (tmp5430 & tmp5434);
  wire tmp5436;
  assign tmp5436 = 1'b0;
  wire tmp5437;
  assign tmp5437 = ~pi7;
  wire tmp5438;
  assign tmp5438 = 1'b0;
  wire tmp5439;
  assign tmp5439 = (tmp5436 & tmp5437) | (tmp5436 & tmp5438) | (tmp5437 & tmp5438);
  wire tmp5440;
  assign tmp5440 = ~pi7;
  wire tmp5441;
  assign tmp5441 = 1'b1;
  wire tmp5442;
  assign tmp5442 = 1'b0;
  wire tmp5443;
  assign tmp5443 = (tmp5440 & tmp5441) | (tmp5440 & tmp5442) | (tmp5441 & tmp5442);
  wire tmp5444;
  assign tmp5444 = 1'b0;
  wire tmp5445;
  assign tmp5445 = 1'b0;
  wire tmp5446;
  assign tmp5446 = 1'b0;
  wire tmp5447;
  assign tmp5447 = (tmp5444 & tmp5445) | (tmp5444 & tmp5446) | (tmp5445 & tmp5446);
  wire tmp5448;
  assign tmp5448 = (tmp5439 & tmp5443) | (tmp5439 & tmp5447) | (tmp5443 & tmp5447);
  wire tmp5449;
  assign tmp5449 = 1'b0;
  wire tmp5450;
  assign tmp5450 = 1'b0;
  wire tmp5451;
  assign tmp5451 = 1'b0;
  wire tmp5452;
  assign tmp5452 = (tmp5449 & tmp5450) | (tmp5449 & tmp5451) | (tmp5450 & tmp5451);
  wire tmp5453;
  assign tmp5453 = 1'b0;
  wire tmp5454;
  assign tmp5454 = 1'b0;
  wire tmp5455;
  assign tmp5455 = 1'b0;
  wire tmp5456;
  assign tmp5456 = (tmp5453 & tmp5454) | (tmp5453 & tmp5455) | (tmp5454 & tmp5455);
  wire tmp5457;
  assign tmp5457 = 1'b0;
  wire tmp5458;
  assign tmp5458 = 1'b0;
  wire tmp5459;
  assign tmp5459 = 1'b0;
  wire tmp5460;
  assign tmp5460 = (tmp5457 & tmp5458) | (tmp5457 & tmp5459) | (tmp5458 & tmp5459);
  wire tmp5461;
  assign tmp5461 = (tmp5452 & tmp5456) | (tmp5452 & tmp5460) | (tmp5456 & tmp5460);
  wire tmp5462;
  assign tmp5462 = (tmp5435 & tmp5448) | (tmp5435 & tmp5461) | (tmp5448 & tmp5461);
  wire tmp5463;
  assign tmp5463 = (tmp5382 & tmp5422) | (tmp5382 & tmp5462) | (tmp5422 & tmp5462);
  wire tmp5464;
  assign tmp5464 = (tmp5221 & tmp5342) | (tmp5221 & tmp5463) | (tmp5342 & tmp5463);
  wire tmp5465;
  assign tmp5465 = (tmp4736 & tmp5100) | (tmp4736 & tmp5464) | (tmp5100 & tmp5464);
  wire tmp5466;
  assign tmp5466 = 1'b0;
  wire tmp5467;
  assign tmp5467 = 1'b0;
  wire tmp5468;
  assign tmp5468 = 1'b0;
  wire tmp5469;
  assign tmp5469 = (tmp5466 & tmp5467) | (tmp5466 & tmp5468) | (tmp5467 & tmp5468);
  wire tmp5470;
  assign tmp5470 = 1'b0;
  wire tmp5471;
  assign tmp5471 = 1'b0;
  wire tmp5472;
  assign tmp5472 = 1'b0;
  wire tmp5473;
  assign tmp5473 = (tmp5470 & tmp5471) | (tmp5470 & tmp5472) | (tmp5471 & tmp5472);
  wire tmp5474;
  assign tmp5474 = 1'b0;
  wire tmp5475;
  assign tmp5475 = 1'b0;
  wire tmp5476;
  assign tmp5476 = 1'b0;
  wire tmp5477;
  assign tmp5477 = (tmp5474 & tmp5475) | (tmp5474 & tmp5476) | (tmp5475 & tmp5476);
  wire tmp5478;
  assign tmp5478 = (tmp5469 & tmp5473) | (tmp5469 & tmp5477) | (tmp5473 & tmp5477);
  wire tmp5479;
  assign tmp5479 = 1'b0;
  wire tmp5480;
  assign tmp5480 = 1'b0;
  wire tmp5481;
  assign tmp5481 = 1'b0;
  wire tmp5482;
  assign tmp5482 = (tmp5479 & tmp5480) | (tmp5479 & tmp5481) | (tmp5480 & tmp5481);
  wire tmp5483;
  assign tmp5483 = 1'b0;
  wire tmp5484;
  assign tmp5484 = 1'b1;
  wire tmp5485;
  assign tmp5485 = 1'b0;
  wire tmp5486;
  assign tmp5486 = (tmp5483 & tmp5484) | (tmp5483 & tmp5485) | (tmp5484 & tmp5485);
  wire tmp5487;
  assign tmp5487 = 1'b0;
  wire tmp5488;
  assign tmp5488 = 1'b0;
  wire tmp5489;
  assign tmp5489 = 1'b0;
  wire tmp5490;
  assign tmp5490 = (tmp5487 & tmp5488) | (tmp5487 & tmp5489) | (tmp5488 & tmp5489);
  wire tmp5491;
  assign tmp5491 = (tmp5482 & tmp5486) | (tmp5482 & tmp5490) | (tmp5486 & tmp5490);
  wire tmp5492;
  assign tmp5492 = 1'b0;
  wire tmp5493;
  assign tmp5493 = 1'b0;
  wire tmp5494;
  assign tmp5494 = 1'b0;
  wire tmp5495;
  assign tmp5495 = (tmp5492 & tmp5493) | (tmp5492 & tmp5494) | (tmp5493 & tmp5494);
  wire tmp5496;
  assign tmp5496 = 1'b0;
  wire tmp5497;
  assign tmp5497 = 1'b0;
  wire tmp5498;
  assign tmp5498 = 1'b0;
  wire tmp5499;
  assign tmp5499 = (tmp5496 & tmp5497) | (tmp5496 & tmp5498) | (tmp5497 & tmp5498);
  wire tmp5500;
  assign tmp5500 = 1'b0;
  wire tmp5501;
  assign tmp5501 = 1'b0;
  wire tmp5502;
  assign tmp5502 = 1'b0;
  wire tmp5503;
  assign tmp5503 = (tmp5500 & tmp5501) | (tmp5500 & tmp5502) | (tmp5501 & tmp5502);
  wire tmp5504;
  assign tmp5504 = (tmp5495 & tmp5499) | (tmp5495 & tmp5503) | (tmp5499 & tmp5503);
  wire tmp5505;
  assign tmp5505 = (tmp5478 & tmp5491) | (tmp5478 & tmp5504) | (tmp5491 & tmp5504);
  wire tmp5506;
  assign tmp5506 = 1'b0;
  wire tmp5507;
  assign tmp5507 = 1'b0;
  wire tmp5508;
  assign tmp5508 = 1'b0;
  wire tmp5509;
  assign tmp5509 = (tmp5506 & tmp5507) | (tmp5506 & tmp5508) | (tmp5507 & tmp5508);
  wire tmp5510;
  assign tmp5510 = 1'b0;
  wire tmp5511;
  assign tmp5511 = 1'b1;
  wire tmp5512;
  assign tmp5512 = 1'b0;
  wire tmp5513;
  assign tmp5513 = (tmp5510 & tmp5511) | (tmp5510 & tmp5512) | (tmp5511 & tmp5512);
  wire tmp5514;
  assign tmp5514 = 1'b0;
  wire tmp5515;
  assign tmp5515 = 1'b0;
  wire tmp5516;
  assign tmp5516 = 1'b0;
  wire tmp5517;
  assign tmp5517 = (tmp5514 & tmp5515) | (tmp5514 & tmp5516) | (tmp5515 & tmp5516);
  wire tmp5518;
  assign tmp5518 = (tmp5509 & tmp5513) | (tmp5509 & tmp5517) | (tmp5513 & tmp5517);
  wire tmp5519;
  assign tmp5519 = 1'b0;
  wire tmp5520;
  assign tmp5520 = 1'b1;
  wire tmp5521;
  assign tmp5521 = 1'b0;
  wire tmp5522;
  assign tmp5522 = (tmp5519 & tmp5520) | (tmp5519 & tmp5521) | (tmp5520 & tmp5521);
  wire tmp5523;
  assign tmp5523 = 1'b1;
  wire tmp5524;
  assign tmp5524 = 1'b1;
  wire tmp5525;
  assign tmp5525 = 1'b1;
  wire tmp5526;
  assign tmp5526 = (tmp5523 & tmp5524) | (tmp5523 & tmp5525) | (tmp5524 & tmp5525);
  wire tmp5527;
  assign tmp5527 = 1'b0;
  wire tmp5528;
  assign tmp5528 = 1'b1;
  wire tmp5529;
  assign tmp5529 = 1'b0;
  wire tmp5530;
  assign tmp5530 = (tmp5527 & tmp5528) | (tmp5527 & tmp5529) | (tmp5528 & tmp5529);
  wire tmp5531;
  assign tmp5531 = (tmp5522 & tmp5526) | (tmp5522 & tmp5530) | (tmp5526 & tmp5530);
  wire tmp5532;
  assign tmp5532 = 1'b0;
  wire tmp5533;
  assign tmp5533 = 1'b0;
  wire tmp5534;
  assign tmp5534 = 1'b0;
  wire tmp5535;
  assign tmp5535 = (tmp5532 & tmp5533) | (tmp5532 & tmp5534) | (tmp5533 & tmp5534);
  wire tmp5536;
  assign tmp5536 = 1'b0;
  wire tmp5537;
  assign tmp5537 = 1'b1;
  wire tmp5538;
  assign tmp5538 = 1'b0;
  wire tmp5539;
  assign tmp5539 = (tmp5536 & tmp5537) | (tmp5536 & tmp5538) | (tmp5537 & tmp5538);
  wire tmp5540;
  assign tmp5540 = 1'b0;
  wire tmp5541;
  assign tmp5541 = 1'b0;
  wire tmp5542;
  assign tmp5542 = 1'b0;
  wire tmp5543;
  assign tmp5543 = (tmp5540 & tmp5541) | (tmp5540 & tmp5542) | (tmp5541 & tmp5542);
  wire tmp5544;
  assign tmp5544 = (tmp5535 & tmp5539) | (tmp5535 & tmp5543) | (tmp5539 & tmp5543);
  wire tmp5545;
  assign tmp5545 = (tmp5518 & tmp5531) | (tmp5518 & tmp5544) | (tmp5531 & tmp5544);
  wire tmp5546;
  assign tmp5546 = 1'b0;
  wire tmp5547;
  assign tmp5547 = 1'b0;
  wire tmp5548;
  assign tmp5548 = 1'b0;
  wire tmp5549;
  assign tmp5549 = (tmp5546 & tmp5547) | (tmp5546 & tmp5548) | (tmp5547 & tmp5548);
  wire tmp5550;
  assign tmp5550 = 1'b0;
  wire tmp5551;
  assign tmp5551 = 1'b0;
  wire tmp5552;
  assign tmp5552 = 1'b0;
  wire tmp5553;
  assign tmp5553 = (tmp5550 & tmp5551) | (tmp5550 & tmp5552) | (tmp5551 & tmp5552);
  wire tmp5554;
  assign tmp5554 = 1'b0;
  wire tmp5555;
  assign tmp5555 = 1'b0;
  wire tmp5556;
  assign tmp5556 = 1'b0;
  wire tmp5557;
  assign tmp5557 = (tmp5554 & tmp5555) | (tmp5554 & tmp5556) | (tmp5555 & tmp5556);
  wire tmp5558;
  assign tmp5558 = (tmp5549 & tmp5553) | (tmp5549 & tmp5557) | (tmp5553 & tmp5557);
  wire tmp5559;
  assign tmp5559 = 1'b0;
  wire tmp5560;
  assign tmp5560 = 1'b0;
  wire tmp5561;
  assign tmp5561 = 1'b0;
  wire tmp5562;
  assign tmp5562 = (tmp5559 & tmp5560) | (tmp5559 & tmp5561) | (tmp5560 & tmp5561);
  wire tmp5563;
  assign tmp5563 = 1'b0;
  wire tmp5564;
  assign tmp5564 = 1'b1;
  wire tmp5565;
  assign tmp5565 = 1'b0;
  wire tmp5566;
  assign tmp5566 = (tmp5563 & tmp5564) | (tmp5563 & tmp5565) | (tmp5564 & tmp5565);
  wire tmp5567;
  assign tmp5567 = 1'b0;
  wire tmp5568;
  assign tmp5568 = 1'b0;
  wire tmp5569;
  assign tmp5569 = 1'b0;
  wire tmp5570;
  assign tmp5570 = (tmp5567 & tmp5568) | (tmp5567 & tmp5569) | (tmp5568 & tmp5569);
  wire tmp5571;
  assign tmp5571 = (tmp5562 & tmp5566) | (tmp5562 & tmp5570) | (tmp5566 & tmp5570);
  wire tmp5572;
  assign tmp5572 = 1'b0;
  wire tmp5573;
  assign tmp5573 = 1'b0;
  wire tmp5574;
  assign tmp5574 = 1'b0;
  wire tmp5575;
  assign tmp5575 = (tmp5572 & tmp5573) | (tmp5572 & tmp5574) | (tmp5573 & tmp5574);
  wire tmp5576;
  assign tmp5576 = 1'b0;
  wire tmp5577;
  assign tmp5577 = 1'b0;
  wire tmp5578;
  assign tmp5578 = 1'b0;
  wire tmp5579;
  assign tmp5579 = (tmp5576 & tmp5577) | (tmp5576 & tmp5578) | (tmp5577 & tmp5578);
  wire tmp5580;
  assign tmp5580 = 1'b0;
  wire tmp5581;
  assign tmp5581 = 1'b0;
  wire tmp5582;
  assign tmp5582 = 1'b0;
  wire tmp5583;
  assign tmp5583 = (tmp5580 & tmp5581) | (tmp5580 & tmp5582) | (tmp5581 & tmp5582);
  wire tmp5584;
  assign tmp5584 = (tmp5575 & tmp5579) | (tmp5575 & tmp5583) | (tmp5579 & tmp5583);
  wire tmp5585;
  assign tmp5585 = (tmp5558 & tmp5571) | (tmp5558 & tmp5584) | (tmp5571 & tmp5584);
  wire tmp5586;
  assign tmp5586 = (tmp5505 & tmp5545) | (tmp5505 & tmp5585) | (tmp5545 & tmp5585);
  wire tmp5587;
  assign tmp5587 = 1'b0;
  wire tmp5588;
  assign tmp5588 = 1'b0;
  wire tmp5589;
  assign tmp5589 = 1'b0;
  wire tmp5590;
  assign tmp5590 = (tmp5587 & tmp5588) | (tmp5587 & tmp5589) | (tmp5588 & tmp5589);
  wire tmp5591;
  assign tmp5591 = 1'b0;
  wire tmp5592;
  assign tmp5592 = 1'b1;
  wire tmp5593;
  assign tmp5593 = 1'b0;
  wire tmp5594;
  assign tmp5594 = (tmp5591 & tmp5592) | (tmp5591 & tmp5593) | (tmp5592 & tmp5593);
  wire tmp5595;
  assign tmp5595 = 1'b0;
  wire tmp5596;
  assign tmp5596 = 1'b0;
  wire tmp5597;
  assign tmp5597 = 1'b0;
  wire tmp5598;
  assign tmp5598 = (tmp5595 & tmp5596) | (tmp5595 & tmp5597) | (tmp5596 & tmp5597);
  wire tmp5599;
  assign tmp5599 = (tmp5590 & tmp5594) | (tmp5590 & tmp5598) | (tmp5594 & tmp5598);
  wire tmp5600;
  assign tmp5600 = 1'b0;
  wire tmp5601;
  assign tmp5601 = 1'b1;
  wire tmp5602;
  assign tmp5602 = 1'b0;
  wire tmp5603;
  assign tmp5603 = (tmp5600 & tmp5601) | (tmp5600 & tmp5602) | (tmp5601 & tmp5602);
  wire tmp5604;
  assign tmp5604 = 1'b1;
  wire tmp5605;
  assign tmp5605 = 1'b1;
  wire tmp5606;
  assign tmp5606 = 1'b1;
  wire tmp5607;
  assign tmp5607 = (tmp5604 & tmp5605) | (tmp5604 & tmp5606) | (tmp5605 & tmp5606);
  wire tmp5608;
  assign tmp5608 = 1'b0;
  wire tmp5609;
  assign tmp5609 = 1'b1;
  wire tmp5610;
  assign tmp5610 = 1'b0;
  wire tmp5611;
  assign tmp5611 = (tmp5608 & tmp5609) | (tmp5608 & tmp5610) | (tmp5609 & tmp5610);
  wire tmp5612;
  assign tmp5612 = (tmp5603 & tmp5607) | (tmp5603 & tmp5611) | (tmp5607 & tmp5611);
  wire tmp5613;
  assign tmp5613 = 1'b0;
  wire tmp5614;
  assign tmp5614 = 1'b0;
  wire tmp5615;
  assign tmp5615 = 1'b0;
  wire tmp5616;
  assign tmp5616 = (tmp5613 & tmp5614) | (tmp5613 & tmp5615) | (tmp5614 & tmp5615);
  wire tmp5617;
  assign tmp5617 = 1'b0;
  wire tmp5618;
  assign tmp5618 = 1'b1;
  wire tmp5619;
  assign tmp5619 = 1'b0;
  wire tmp5620;
  assign tmp5620 = (tmp5617 & tmp5618) | (tmp5617 & tmp5619) | (tmp5618 & tmp5619);
  wire tmp5621;
  assign tmp5621 = 1'b0;
  wire tmp5622;
  assign tmp5622 = 1'b0;
  wire tmp5623;
  assign tmp5623 = 1'b0;
  wire tmp5624;
  assign tmp5624 = (tmp5621 & tmp5622) | (tmp5621 & tmp5623) | (tmp5622 & tmp5623);
  wire tmp5625;
  assign tmp5625 = (tmp5616 & tmp5620) | (tmp5616 & tmp5624) | (tmp5620 & tmp5624);
  wire tmp5626;
  assign tmp5626 = (tmp5599 & tmp5612) | (tmp5599 & tmp5625) | (tmp5612 & tmp5625);
  wire tmp5627;
  assign tmp5627 = 1'b0;
  wire tmp5628;
  assign tmp5628 = 1'b1;
  wire tmp5629;
  assign tmp5629 = 1'b0;
  wire tmp5630;
  assign tmp5630 = (tmp5627 & tmp5628) | (tmp5627 & tmp5629) | (tmp5628 & tmp5629);
  wire tmp5631;
  assign tmp5631 = 1'b1;
  wire tmp5632;
  assign tmp5632 = 1'b1;
  wire tmp5633;
  assign tmp5633 = 1'b1;
  wire tmp5634;
  assign tmp5634 = (tmp5631 & tmp5632) | (tmp5631 & tmp5633) | (tmp5632 & tmp5633);
  wire tmp5635;
  assign tmp5635 = 1'b0;
  wire tmp5636;
  assign tmp5636 = 1'b1;
  wire tmp5637;
  assign tmp5637 = 1'b0;
  wire tmp5638;
  assign tmp5638 = (tmp5635 & tmp5636) | (tmp5635 & tmp5637) | (tmp5636 & tmp5637);
  wire tmp5639;
  assign tmp5639 = (tmp5630 & tmp5634) | (tmp5630 & tmp5638) | (tmp5634 & tmp5638);
  wire tmp5640;
  assign tmp5640 = 1'b1;
  wire tmp5641;
  assign tmp5641 = 1'b1;
  wire tmp5642;
  assign tmp5642 = 1'b1;
  wire tmp5643;
  assign tmp5643 = (tmp5640 & tmp5641) | (tmp5640 & tmp5642) | (tmp5641 & tmp5642);
  wire tmp5644;
  assign tmp5644 = 1'b1;
  wire tmp5645;
  assign tmp5645 = ~pi5;
  wire tmp5646;
  assign tmp5646 = ~pi6;
  wire tmp5647;
  assign tmp5647 = (tmp5644 & tmp5645) | (tmp5644 & tmp5646) | (tmp5645 & tmp5646);
  wire tmp5648;
  assign tmp5648 = 1'b1;
  wire tmp5649;
  assign tmp5649 = ~pi6;
  wire tmp5650;
  assign tmp5650 = ~pi7;
  wire tmp5651;
  assign tmp5651 = (tmp5648 & tmp5649) | (tmp5648 & tmp5650) | (tmp5649 & tmp5650);
  wire tmp5652;
  assign tmp5652 = (tmp5643 & tmp5647) | (tmp5643 & tmp5651) | (tmp5647 & tmp5651);
  wire tmp5653;
  assign tmp5653 = 1'b0;
  wire tmp5654;
  assign tmp5654 = 1'b1;
  wire tmp5655;
  assign tmp5655 = 1'b0;
  wire tmp5656;
  assign tmp5656 = (tmp5653 & tmp5654) | (tmp5653 & tmp5655) | (tmp5654 & tmp5655);
  wire tmp5657;
  assign tmp5657 = 1'b1;
  wire tmp5658;
  assign tmp5658 = ~pi6;
  wire tmp5659;
  assign tmp5659 = ~pi7;
  wire tmp5660;
  assign tmp5660 = (tmp5657 & tmp5658) | (tmp5657 & tmp5659) | (tmp5658 & tmp5659);
  wire tmp5661;
  assign tmp5661 = 1'b0;
  wire tmp5662;
  assign tmp5662 = ~pi7;
  wire tmp5663;
  assign tmp5663 = 1'b0;
  wire tmp5664;
  assign tmp5664 = (tmp5661 & tmp5662) | (tmp5661 & tmp5663) | (tmp5662 & tmp5663);
  wire tmp5665;
  assign tmp5665 = (tmp5656 & tmp5660) | (tmp5656 & tmp5664) | (tmp5660 & tmp5664);
  wire tmp5666;
  assign tmp5666 = (tmp5639 & tmp5652) | (tmp5639 & tmp5665) | (tmp5652 & tmp5665);
  wire tmp5667;
  assign tmp5667 = 1'b0;
  wire tmp5668;
  assign tmp5668 = 1'b0;
  wire tmp5669;
  assign tmp5669 = 1'b0;
  wire tmp5670;
  assign tmp5670 = (tmp5667 & tmp5668) | (tmp5667 & tmp5669) | (tmp5668 & tmp5669);
  wire tmp5671;
  assign tmp5671 = 1'b0;
  wire tmp5672;
  assign tmp5672 = 1'b1;
  wire tmp5673;
  assign tmp5673 = 1'b0;
  wire tmp5674;
  assign tmp5674 = (tmp5671 & tmp5672) | (tmp5671 & tmp5673) | (tmp5672 & tmp5673);
  wire tmp5675;
  assign tmp5675 = 1'b0;
  wire tmp5676;
  assign tmp5676 = 1'b0;
  wire tmp5677;
  assign tmp5677 = 1'b0;
  wire tmp5678;
  assign tmp5678 = (tmp5675 & tmp5676) | (tmp5675 & tmp5677) | (tmp5676 & tmp5677);
  wire tmp5679;
  assign tmp5679 = (tmp5670 & tmp5674) | (tmp5670 & tmp5678) | (tmp5674 & tmp5678);
  wire tmp5680;
  assign tmp5680 = 1'b0;
  wire tmp5681;
  assign tmp5681 = 1'b1;
  wire tmp5682;
  assign tmp5682 = 1'b0;
  wire tmp5683;
  assign tmp5683 = (tmp5680 & tmp5681) | (tmp5680 & tmp5682) | (tmp5681 & tmp5682);
  wire tmp5684;
  assign tmp5684 = 1'b1;
  wire tmp5685;
  assign tmp5685 = ~pi6;
  wire tmp5686;
  assign tmp5686 = ~pi7;
  wire tmp5687;
  assign tmp5687 = (tmp5684 & tmp5685) | (tmp5684 & tmp5686) | (tmp5685 & tmp5686);
  wire tmp5688;
  assign tmp5688 = 1'b0;
  wire tmp5689;
  assign tmp5689 = ~pi7;
  wire tmp5690;
  assign tmp5690 = 1'b0;
  wire tmp5691;
  assign tmp5691 = (tmp5688 & tmp5689) | (tmp5688 & tmp5690) | (tmp5689 & tmp5690);
  wire tmp5692;
  assign tmp5692 = (tmp5683 & tmp5687) | (tmp5683 & tmp5691) | (tmp5687 & tmp5691);
  wire tmp5693;
  assign tmp5693 = 1'b0;
  wire tmp5694;
  assign tmp5694 = 1'b0;
  wire tmp5695;
  assign tmp5695 = 1'b0;
  wire tmp5696;
  assign tmp5696 = (tmp5693 & tmp5694) | (tmp5693 & tmp5695) | (tmp5694 & tmp5695);
  wire tmp5697;
  assign tmp5697 = 1'b0;
  wire tmp5698;
  assign tmp5698 = ~pi7;
  wire tmp5699;
  assign tmp5699 = 1'b0;
  wire tmp5700;
  assign tmp5700 = (tmp5697 & tmp5698) | (tmp5697 & tmp5699) | (tmp5698 & tmp5699);
  wire tmp5701;
  assign tmp5701 = 1'b0;
  wire tmp5702;
  assign tmp5702 = 1'b0;
  wire tmp5703;
  assign tmp5703 = 1'b0;
  wire tmp5704;
  assign tmp5704 = (tmp5701 & tmp5702) | (tmp5701 & tmp5703) | (tmp5702 & tmp5703);
  wire tmp5705;
  assign tmp5705 = (tmp5696 & tmp5700) | (tmp5696 & tmp5704) | (tmp5700 & tmp5704);
  wire tmp5706;
  assign tmp5706 = (tmp5679 & tmp5692) | (tmp5679 & tmp5705) | (tmp5692 & tmp5705);
  wire tmp5707;
  assign tmp5707 = (tmp5626 & tmp5666) | (tmp5626 & tmp5706) | (tmp5666 & tmp5706);
  wire tmp5708;
  assign tmp5708 = 1'b0;
  wire tmp5709;
  assign tmp5709 = 1'b0;
  wire tmp5710;
  assign tmp5710 = 1'b0;
  wire tmp5711;
  assign tmp5711 = (tmp5708 & tmp5709) | (tmp5708 & tmp5710) | (tmp5709 & tmp5710);
  wire tmp5712;
  assign tmp5712 = 1'b0;
  wire tmp5713;
  assign tmp5713 = 1'b0;
  wire tmp5714;
  assign tmp5714 = 1'b0;
  wire tmp5715;
  assign tmp5715 = (tmp5712 & tmp5713) | (tmp5712 & tmp5714) | (tmp5713 & tmp5714);
  wire tmp5716;
  assign tmp5716 = 1'b0;
  wire tmp5717;
  assign tmp5717 = 1'b0;
  wire tmp5718;
  assign tmp5718 = 1'b0;
  wire tmp5719;
  assign tmp5719 = (tmp5716 & tmp5717) | (tmp5716 & tmp5718) | (tmp5717 & tmp5718);
  wire tmp5720;
  assign tmp5720 = (tmp5711 & tmp5715) | (tmp5711 & tmp5719) | (tmp5715 & tmp5719);
  wire tmp5721;
  assign tmp5721 = 1'b0;
  wire tmp5722;
  assign tmp5722 = 1'b0;
  wire tmp5723;
  assign tmp5723 = 1'b0;
  wire tmp5724;
  assign tmp5724 = (tmp5721 & tmp5722) | (tmp5721 & tmp5723) | (tmp5722 & tmp5723);
  wire tmp5725;
  assign tmp5725 = 1'b0;
  wire tmp5726;
  assign tmp5726 = 1'b1;
  wire tmp5727;
  assign tmp5727 = 1'b0;
  wire tmp5728;
  assign tmp5728 = (tmp5725 & tmp5726) | (tmp5725 & tmp5727) | (tmp5726 & tmp5727);
  wire tmp5729;
  assign tmp5729 = 1'b0;
  wire tmp5730;
  assign tmp5730 = 1'b0;
  wire tmp5731;
  assign tmp5731 = 1'b0;
  wire tmp5732;
  assign tmp5732 = (tmp5729 & tmp5730) | (tmp5729 & tmp5731) | (tmp5730 & tmp5731);
  wire tmp5733;
  assign tmp5733 = (tmp5724 & tmp5728) | (tmp5724 & tmp5732) | (tmp5728 & tmp5732);
  wire tmp5734;
  assign tmp5734 = 1'b0;
  wire tmp5735;
  assign tmp5735 = 1'b0;
  wire tmp5736;
  assign tmp5736 = 1'b0;
  wire tmp5737;
  assign tmp5737 = (tmp5734 & tmp5735) | (tmp5734 & tmp5736) | (tmp5735 & tmp5736);
  wire tmp5738;
  assign tmp5738 = 1'b0;
  wire tmp5739;
  assign tmp5739 = 1'b0;
  wire tmp5740;
  assign tmp5740 = 1'b0;
  wire tmp5741;
  assign tmp5741 = (tmp5738 & tmp5739) | (tmp5738 & tmp5740) | (tmp5739 & tmp5740);
  wire tmp5742;
  assign tmp5742 = 1'b0;
  wire tmp5743;
  assign tmp5743 = 1'b0;
  wire tmp5744;
  assign tmp5744 = 1'b0;
  wire tmp5745;
  assign tmp5745 = (tmp5742 & tmp5743) | (tmp5742 & tmp5744) | (tmp5743 & tmp5744);
  wire tmp5746;
  assign tmp5746 = (tmp5737 & tmp5741) | (tmp5737 & tmp5745) | (tmp5741 & tmp5745);
  wire tmp5747;
  assign tmp5747 = (tmp5720 & tmp5733) | (tmp5720 & tmp5746) | (tmp5733 & tmp5746);
  wire tmp5748;
  assign tmp5748 = 1'b0;
  wire tmp5749;
  assign tmp5749 = 1'b0;
  wire tmp5750;
  assign tmp5750 = 1'b0;
  wire tmp5751;
  assign tmp5751 = (tmp5748 & tmp5749) | (tmp5748 & tmp5750) | (tmp5749 & tmp5750);
  wire tmp5752;
  assign tmp5752 = 1'b0;
  wire tmp5753;
  assign tmp5753 = 1'b1;
  wire tmp5754;
  assign tmp5754 = 1'b0;
  wire tmp5755;
  assign tmp5755 = (tmp5752 & tmp5753) | (tmp5752 & tmp5754) | (tmp5753 & tmp5754);
  wire tmp5756;
  assign tmp5756 = 1'b0;
  wire tmp5757;
  assign tmp5757 = 1'b0;
  wire tmp5758;
  assign tmp5758 = 1'b0;
  wire tmp5759;
  assign tmp5759 = (tmp5756 & tmp5757) | (tmp5756 & tmp5758) | (tmp5757 & tmp5758);
  wire tmp5760;
  assign tmp5760 = (tmp5751 & tmp5755) | (tmp5751 & tmp5759) | (tmp5755 & tmp5759);
  wire tmp5761;
  assign tmp5761 = 1'b0;
  wire tmp5762;
  assign tmp5762 = 1'b1;
  wire tmp5763;
  assign tmp5763 = 1'b0;
  wire tmp5764;
  assign tmp5764 = (tmp5761 & tmp5762) | (tmp5761 & tmp5763) | (tmp5762 & tmp5763);
  wire tmp5765;
  assign tmp5765 = 1'b1;
  wire tmp5766;
  assign tmp5766 = ~pi6;
  wire tmp5767;
  assign tmp5767 = ~pi7;
  wire tmp5768;
  assign tmp5768 = (tmp5765 & tmp5766) | (tmp5765 & tmp5767) | (tmp5766 & tmp5767);
  wire tmp5769;
  assign tmp5769 = 1'b0;
  wire tmp5770;
  assign tmp5770 = ~pi7;
  wire tmp5771;
  assign tmp5771 = 1'b0;
  wire tmp5772;
  assign tmp5772 = (tmp5769 & tmp5770) | (tmp5769 & tmp5771) | (tmp5770 & tmp5771);
  wire tmp5773;
  assign tmp5773 = (tmp5764 & tmp5768) | (tmp5764 & tmp5772) | (tmp5768 & tmp5772);
  wire tmp5774;
  assign tmp5774 = 1'b0;
  wire tmp5775;
  assign tmp5775 = 1'b0;
  wire tmp5776;
  assign tmp5776 = 1'b0;
  wire tmp5777;
  assign tmp5777 = (tmp5774 & tmp5775) | (tmp5774 & tmp5776) | (tmp5775 & tmp5776);
  wire tmp5778;
  assign tmp5778 = 1'b0;
  wire tmp5779;
  assign tmp5779 = ~pi7;
  wire tmp5780;
  assign tmp5780 = 1'b0;
  wire tmp5781;
  assign tmp5781 = (tmp5778 & tmp5779) | (tmp5778 & tmp5780) | (tmp5779 & tmp5780);
  wire tmp5782;
  assign tmp5782 = 1'b0;
  wire tmp5783;
  assign tmp5783 = 1'b0;
  wire tmp5784;
  assign tmp5784 = 1'b0;
  wire tmp5785;
  assign tmp5785 = (tmp5782 & tmp5783) | (tmp5782 & tmp5784) | (tmp5783 & tmp5784);
  wire tmp5786;
  assign tmp5786 = (tmp5777 & tmp5781) | (tmp5777 & tmp5785) | (tmp5781 & tmp5785);
  wire tmp5787;
  assign tmp5787 = (tmp5760 & tmp5773) | (tmp5760 & tmp5786) | (tmp5773 & tmp5786);
  wire tmp5788;
  assign tmp5788 = 1'b0;
  wire tmp5789;
  assign tmp5789 = 1'b0;
  wire tmp5790;
  assign tmp5790 = 1'b0;
  wire tmp5791;
  assign tmp5791 = (tmp5788 & tmp5789) | (tmp5788 & tmp5790) | (tmp5789 & tmp5790);
  wire tmp5792;
  assign tmp5792 = 1'b0;
  wire tmp5793;
  assign tmp5793 = 1'b0;
  wire tmp5794;
  assign tmp5794 = 1'b0;
  wire tmp5795;
  assign tmp5795 = (tmp5792 & tmp5793) | (tmp5792 & tmp5794) | (tmp5793 & tmp5794);
  wire tmp5796;
  assign tmp5796 = 1'b0;
  wire tmp5797;
  assign tmp5797 = 1'b0;
  wire tmp5798;
  assign tmp5798 = 1'b0;
  wire tmp5799;
  assign tmp5799 = (tmp5796 & tmp5797) | (tmp5796 & tmp5798) | (tmp5797 & tmp5798);
  wire tmp5800;
  assign tmp5800 = (tmp5791 & tmp5795) | (tmp5791 & tmp5799) | (tmp5795 & tmp5799);
  wire tmp5801;
  assign tmp5801 = 1'b0;
  wire tmp5802;
  assign tmp5802 = 1'b0;
  wire tmp5803;
  assign tmp5803 = 1'b0;
  wire tmp5804;
  assign tmp5804 = (tmp5801 & tmp5802) | (tmp5801 & tmp5803) | (tmp5802 & tmp5803);
  wire tmp5805;
  assign tmp5805 = 1'b0;
  wire tmp5806;
  assign tmp5806 = ~pi7;
  wire tmp5807;
  assign tmp5807 = 1'b0;
  wire tmp5808;
  assign tmp5808 = (tmp5805 & tmp5806) | (tmp5805 & tmp5807) | (tmp5806 & tmp5807);
  wire tmp5809;
  assign tmp5809 = 1'b0;
  wire tmp5810;
  assign tmp5810 = 1'b0;
  wire tmp5811;
  assign tmp5811 = 1'b0;
  wire tmp5812;
  assign tmp5812 = (tmp5809 & tmp5810) | (tmp5809 & tmp5811) | (tmp5810 & tmp5811);
  wire tmp5813;
  assign tmp5813 = (tmp5804 & tmp5808) | (tmp5804 & tmp5812) | (tmp5808 & tmp5812);
  wire tmp5814;
  assign tmp5814 = 1'b0;
  wire tmp5815;
  assign tmp5815 = 1'b0;
  wire tmp5816;
  assign tmp5816 = 1'b0;
  wire tmp5817;
  assign tmp5817 = (tmp5814 & tmp5815) | (tmp5814 & tmp5816) | (tmp5815 & tmp5816);
  wire tmp5818;
  assign tmp5818 = 1'b0;
  wire tmp5819;
  assign tmp5819 = 1'b0;
  wire tmp5820;
  assign tmp5820 = 1'b0;
  wire tmp5821;
  assign tmp5821 = (tmp5818 & tmp5819) | (tmp5818 & tmp5820) | (tmp5819 & tmp5820);
  wire tmp5822;
  assign tmp5822 = 1'b0;
  wire tmp5823;
  assign tmp5823 = 1'b0;
  wire tmp5824;
  assign tmp5824 = 1'b0;
  wire tmp5825;
  assign tmp5825 = (tmp5822 & tmp5823) | (tmp5822 & tmp5824) | (tmp5823 & tmp5824);
  wire tmp5826;
  assign tmp5826 = (tmp5817 & tmp5821) | (tmp5817 & tmp5825) | (tmp5821 & tmp5825);
  wire tmp5827;
  assign tmp5827 = (tmp5800 & tmp5813) | (tmp5800 & tmp5826) | (tmp5813 & tmp5826);
  wire tmp5828;
  assign tmp5828 = (tmp5747 & tmp5787) | (tmp5747 & tmp5827) | (tmp5787 & tmp5827);
  wire tmp5829;
  assign tmp5829 = (tmp5586 & tmp5707) | (tmp5586 & tmp5828) | (tmp5707 & tmp5828);
  wire tmp5830;
  assign tmp5830 = 1'b0;
  wire tmp5831;
  assign tmp5831 = 1'b0;
  wire tmp5832;
  assign tmp5832 = 1'b0;
  wire tmp5833;
  assign tmp5833 = (tmp5830 & tmp5831) | (tmp5830 & tmp5832) | (tmp5831 & tmp5832);
  wire tmp5834;
  assign tmp5834 = 1'b0;
  wire tmp5835;
  assign tmp5835 = 1'b1;
  wire tmp5836;
  assign tmp5836 = 1'b0;
  wire tmp5837;
  assign tmp5837 = (tmp5834 & tmp5835) | (tmp5834 & tmp5836) | (tmp5835 & tmp5836);
  wire tmp5838;
  assign tmp5838 = 1'b0;
  wire tmp5839;
  assign tmp5839 = 1'b0;
  wire tmp5840;
  assign tmp5840 = 1'b0;
  wire tmp5841;
  assign tmp5841 = (tmp5838 & tmp5839) | (tmp5838 & tmp5840) | (tmp5839 & tmp5840);
  wire tmp5842;
  assign tmp5842 = (tmp5833 & tmp5837) | (tmp5833 & tmp5841) | (tmp5837 & tmp5841);
  wire tmp5843;
  assign tmp5843 = 1'b0;
  wire tmp5844;
  assign tmp5844 = 1'b1;
  wire tmp5845;
  assign tmp5845 = 1'b0;
  wire tmp5846;
  assign tmp5846 = (tmp5843 & tmp5844) | (tmp5843 & tmp5845) | (tmp5844 & tmp5845);
  wire tmp5847;
  assign tmp5847 = 1'b1;
  wire tmp5848;
  assign tmp5848 = 1'b1;
  wire tmp5849;
  assign tmp5849 = 1'b1;
  wire tmp5850;
  assign tmp5850 = (tmp5847 & tmp5848) | (tmp5847 & tmp5849) | (tmp5848 & tmp5849);
  wire tmp5851;
  assign tmp5851 = 1'b0;
  wire tmp5852;
  assign tmp5852 = 1'b1;
  wire tmp5853;
  assign tmp5853 = 1'b0;
  wire tmp5854;
  assign tmp5854 = (tmp5851 & tmp5852) | (tmp5851 & tmp5853) | (tmp5852 & tmp5853);
  wire tmp5855;
  assign tmp5855 = (tmp5846 & tmp5850) | (tmp5846 & tmp5854) | (tmp5850 & tmp5854);
  wire tmp5856;
  assign tmp5856 = 1'b0;
  wire tmp5857;
  assign tmp5857 = 1'b0;
  wire tmp5858;
  assign tmp5858 = 1'b0;
  wire tmp5859;
  assign tmp5859 = (tmp5856 & tmp5857) | (tmp5856 & tmp5858) | (tmp5857 & tmp5858);
  wire tmp5860;
  assign tmp5860 = 1'b0;
  wire tmp5861;
  assign tmp5861 = 1'b1;
  wire tmp5862;
  assign tmp5862 = 1'b0;
  wire tmp5863;
  assign tmp5863 = (tmp5860 & tmp5861) | (tmp5860 & tmp5862) | (tmp5861 & tmp5862);
  wire tmp5864;
  assign tmp5864 = 1'b0;
  wire tmp5865;
  assign tmp5865 = 1'b0;
  wire tmp5866;
  assign tmp5866 = 1'b0;
  wire tmp5867;
  assign tmp5867 = (tmp5864 & tmp5865) | (tmp5864 & tmp5866) | (tmp5865 & tmp5866);
  wire tmp5868;
  assign tmp5868 = (tmp5859 & tmp5863) | (tmp5859 & tmp5867) | (tmp5863 & tmp5867);
  wire tmp5869;
  assign tmp5869 = (tmp5842 & tmp5855) | (tmp5842 & tmp5868) | (tmp5855 & tmp5868);
  wire tmp5870;
  assign tmp5870 = 1'b0;
  wire tmp5871;
  assign tmp5871 = 1'b1;
  wire tmp5872;
  assign tmp5872 = 1'b0;
  wire tmp5873;
  assign tmp5873 = (tmp5870 & tmp5871) | (tmp5870 & tmp5872) | (tmp5871 & tmp5872);
  wire tmp5874;
  assign tmp5874 = 1'b1;
  wire tmp5875;
  assign tmp5875 = 1'b1;
  wire tmp5876;
  assign tmp5876 = 1'b1;
  wire tmp5877;
  assign tmp5877 = (tmp5874 & tmp5875) | (tmp5874 & tmp5876) | (tmp5875 & tmp5876);
  wire tmp5878;
  assign tmp5878 = 1'b0;
  wire tmp5879;
  assign tmp5879 = 1'b1;
  wire tmp5880;
  assign tmp5880 = 1'b0;
  wire tmp5881;
  assign tmp5881 = (tmp5878 & tmp5879) | (tmp5878 & tmp5880) | (tmp5879 & tmp5880);
  wire tmp5882;
  assign tmp5882 = (tmp5873 & tmp5877) | (tmp5873 & tmp5881) | (tmp5877 & tmp5881);
  wire tmp5883;
  assign tmp5883 = 1'b1;
  wire tmp5884;
  assign tmp5884 = 1'b1;
  wire tmp5885;
  assign tmp5885 = 1'b1;
  wire tmp5886;
  assign tmp5886 = (tmp5883 & tmp5884) | (tmp5883 & tmp5885) | (tmp5884 & tmp5885);
  wire tmp5887;
  assign tmp5887 = 1'b1;
  wire tmp5888;
  assign tmp5888 = ~pi5;
  wire tmp5889;
  assign tmp5889 = ~pi6;
  wire tmp5890;
  assign tmp5890 = (tmp5887 & tmp5888) | (tmp5887 & tmp5889) | (tmp5888 & tmp5889);
  wire tmp5891;
  assign tmp5891 = 1'b1;
  wire tmp5892;
  assign tmp5892 = ~pi6;
  wire tmp5893;
  assign tmp5893 = ~pi7;
  wire tmp5894;
  assign tmp5894 = (tmp5891 & tmp5892) | (tmp5891 & tmp5893) | (tmp5892 & tmp5893);
  wire tmp5895;
  assign tmp5895 = (tmp5886 & tmp5890) | (tmp5886 & tmp5894) | (tmp5890 & tmp5894);
  wire tmp5896;
  assign tmp5896 = 1'b0;
  wire tmp5897;
  assign tmp5897 = 1'b1;
  wire tmp5898;
  assign tmp5898 = 1'b0;
  wire tmp5899;
  assign tmp5899 = (tmp5896 & tmp5897) | (tmp5896 & tmp5898) | (tmp5897 & tmp5898);
  wire tmp5900;
  assign tmp5900 = 1'b1;
  wire tmp5901;
  assign tmp5901 = ~pi6;
  wire tmp5902;
  assign tmp5902 = ~pi7;
  wire tmp5903;
  assign tmp5903 = (tmp5900 & tmp5901) | (tmp5900 & tmp5902) | (tmp5901 & tmp5902);
  wire tmp5904;
  assign tmp5904 = 1'b0;
  wire tmp5905;
  assign tmp5905 = ~pi7;
  wire tmp5906;
  assign tmp5906 = 1'b0;
  wire tmp5907;
  assign tmp5907 = (tmp5904 & tmp5905) | (tmp5904 & tmp5906) | (tmp5905 & tmp5906);
  wire tmp5908;
  assign tmp5908 = (tmp5899 & tmp5903) | (tmp5899 & tmp5907) | (tmp5903 & tmp5907);
  wire tmp5909;
  assign tmp5909 = (tmp5882 & tmp5895) | (tmp5882 & tmp5908) | (tmp5895 & tmp5908);
  wire tmp5910;
  assign tmp5910 = 1'b0;
  wire tmp5911;
  assign tmp5911 = 1'b0;
  wire tmp5912;
  assign tmp5912 = 1'b0;
  wire tmp5913;
  assign tmp5913 = (tmp5910 & tmp5911) | (tmp5910 & tmp5912) | (tmp5911 & tmp5912);
  wire tmp5914;
  assign tmp5914 = 1'b0;
  wire tmp5915;
  assign tmp5915 = 1'b1;
  wire tmp5916;
  assign tmp5916 = 1'b0;
  wire tmp5917;
  assign tmp5917 = (tmp5914 & tmp5915) | (tmp5914 & tmp5916) | (tmp5915 & tmp5916);
  wire tmp5918;
  assign tmp5918 = 1'b0;
  wire tmp5919;
  assign tmp5919 = 1'b0;
  wire tmp5920;
  assign tmp5920 = 1'b0;
  wire tmp5921;
  assign tmp5921 = (tmp5918 & tmp5919) | (tmp5918 & tmp5920) | (tmp5919 & tmp5920);
  wire tmp5922;
  assign tmp5922 = (tmp5913 & tmp5917) | (tmp5913 & tmp5921) | (tmp5917 & tmp5921);
  wire tmp5923;
  assign tmp5923 = 1'b0;
  wire tmp5924;
  assign tmp5924 = 1'b1;
  wire tmp5925;
  assign tmp5925 = 1'b0;
  wire tmp5926;
  assign tmp5926 = (tmp5923 & tmp5924) | (tmp5923 & tmp5925) | (tmp5924 & tmp5925);
  wire tmp5927;
  assign tmp5927 = 1'b1;
  wire tmp5928;
  assign tmp5928 = ~pi6;
  wire tmp5929;
  assign tmp5929 = ~pi7;
  wire tmp5930;
  assign tmp5930 = (tmp5927 & tmp5928) | (tmp5927 & tmp5929) | (tmp5928 & tmp5929);
  wire tmp5931;
  assign tmp5931 = 1'b0;
  wire tmp5932;
  assign tmp5932 = ~pi7;
  wire tmp5933;
  assign tmp5933 = 1'b0;
  wire tmp5934;
  assign tmp5934 = (tmp5931 & tmp5932) | (tmp5931 & tmp5933) | (tmp5932 & tmp5933);
  wire tmp5935;
  assign tmp5935 = (tmp5926 & tmp5930) | (tmp5926 & tmp5934) | (tmp5930 & tmp5934);
  wire tmp5936;
  assign tmp5936 = 1'b0;
  wire tmp5937;
  assign tmp5937 = 1'b0;
  wire tmp5938;
  assign tmp5938 = 1'b0;
  wire tmp5939;
  assign tmp5939 = (tmp5936 & tmp5937) | (tmp5936 & tmp5938) | (tmp5937 & tmp5938);
  wire tmp5940;
  assign tmp5940 = 1'b0;
  wire tmp5941;
  assign tmp5941 = ~pi7;
  wire tmp5942;
  assign tmp5942 = 1'b0;
  wire tmp5943;
  assign tmp5943 = (tmp5940 & tmp5941) | (tmp5940 & tmp5942) | (tmp5941 & tmp5942);
  wire tmp5944;
  assign tmp5944 = 1'b0;
  wire tmp5945;
  assign tmp5945 = 1'b0;
  wire tmp5946;
  assign tmp5946 = 1'b0;
  wire tmp5947;
  assign tmp5947 = (tmp5944 & tmp5945) | (tmp5944 & tmp5946) | (tmp5945 & tmp5946);
  wire tmp5948;
  assign tmp5948 = (tmp5939 & tmp5943) | (tmp5939 & tmp5947) | (tmp5943 & tmp5947);
  wire tmp5949;
  assign tmp5949 = (tmp5922 & tmp5935) | (tmp5922 & tmp5948) | (tmp5935 & tmp5948);
  wire tmp5950;
  assign tmp5950 = (tmp5869 & tmp5909) | (tmp5869 & tmp5949) | (tmp5909 & tmp5949);
  wire tmp5951;
  assign tmp5951 = 1'b0;
  wire tmp5952;
  assign tmp5952 = 1'b1;
  wire tmp5953;
  assign tmp5953 = 1'b0;
  wire tmp5954;
  assign tmp5954 = (tmp5951 & tmp5952) | (tmp5951 & tmp5953) | (tmp5952 & tmp5953);
  wire tmp5955;
  assign tmp5955 = 1'b1;
  wire tmp5956;
  assign tmp5956 = 1'b1;
  wire tmp5957;
  assign tmp5957 = 1'b1;
  wire tmp5958;
  assign tmp5958 = (tmp5955 & tmp5956) | (tmp5955 & tmp5957) | (tmp5956 & tmp5957);
  wire tmp5959;
  assign tmp5959 = 1'b0;
  wire tmp5960;
  assign tmp5960 = 1'b1;
  wire tmp5961;
  assign tmp5961 = 1'b0;
  wire tmp5962;
  assign tmp5962 = (tmp5959 & tmp5960) | (tmp5959 & tmp5961) | (tmp5960 & tmp5961);
  wire tmp5963;
  assign tmp5963 = (tmp5954 & tmp5958) | (tmp5954 & tmp5962) | (tmp5958 & tmp5962);
  wire tmp5964;
  assign tmp5964 = 1'b1;
  wire tmp5965;
  assign tmp5965 = 1'b1;
  wire tmp5966;
  assign tmp5966 = 1'b1;
  wire tmp5967;
  assign tmp5967 = (tmp5964 & tmp5965) | (tmp5964 & tmp5966) | (tmp5965 & tmp5966);
  wire tmp5968;
  assign tmp5968 = 1'b1;
  wire tmp5969;
  assign tmp5969 = ~pi5;
  wire tmp5970;
  assign tmp5970 = ~pi6;
  wire tmp5971;
  assign tmp5971 = (tmp5968 & tmp5969) | (tmp5968 & tmp5970) | (tmp5969 & tmp5970);
  wire tmp5972;
  assign tmp5972 = 1'b1;
  wire tmp5973;
  assign tmp5973 = ~pi6;
  wire tmp5974;
  assign tmp5974 = ~pi7;
  wire tmp5975;
  assign tmp5975 = (tmp5972 & tmp5973) | (tmp5972 & tmp5974) | (tmp5973 & tmp5974);
  wire tmp5976;
  assign tmp5976 = (tmp5967 & tmp5971) | (tmp5967 & tmp5975) | (tmp5971 & tmp5975);
  wire tmp5977;
  assign tmp5977 = 1'b0;
  wire tmp5978;
  assign tmp5978 = 1'b1;
  wire tmp5979;
  assign tmp5979 = 1'b0;
  wire tmp5980;
  assign tmp5980 = (tmp5977 & tmp5978) | (tmp5977 & tmp5979) | (tmp5978 & tmp5979);
  wire tmp5981;
  assign tmp5981 = 1'b1;
  wire tmp5982;
  assign tmp5982 = ~pi6;
  wire tmp5983;
  assign tmp5983 = ~pi7;
  wire tmp5984;
  assign tmp5984 = (tmp5981 & tmp5982) | (tmp5981 & tmp5983) | (tmp5982 & tmp5983);
  wire tmp5985;
  assign tmp5985 = 1'b0;
  wire tmp5986;
  assign tmp5986 = ~pi7;
  wire tmp5987;
  assign tmp5987 = 1'b0;
  wire tmp5988;
  assign tmp5988 = (tmp5985 & tmp5986) | (tmp5985 & tmp5987) | (tmp5986 & tmp5987);
  wire tmp5989;
  assign tmp5989 = (tmp5980 & tmp5984) | (tmp5980 & tmp5988) | (tmp5984 & tmp5988);
  wire tmp5990;
  assign tmp5990 = (tmp5963 & tmp5976) | (tmp5963 & tmp5989) | (tmp5976 & tmp5989);
  wire tmp5991;
  assign tmp5991 = 1'b1;
  wire tmp5992;
  assign tmp5992 = 1'b1;
  wire tmp5993;
  assign tmp5993 = 1'b1;
  wire tmp5994;
  assign tmp5994 = (tmp5991 & tmp5992) | (tmp5991 & tmp5993) | (tmp5992 & tmp5993);
  wire tmp5995;
  assign tmp5995 = 1'b1;
  wire tmp5996;
  assign tmp5996 = ~pi5;
  wire tmp5997;
  assign tmp5997 = ~pi6;
  wire tmp5998;
  assign tmp5998 = (tmp5995 & tmp5996) | (tmp5995 & tmp5997) | (tmp5996 & tmp5997);
  wire tmp5999;
  assign tmp5999 = 1'b1;
  wire tmp6000;
  assign tmp6000 = ~pi6;
  wire tmp6001;
  assign tmp6001 = ~pi7;
  wire tmp6002;
  assign tmp6002 = (tmp5999 & tmp6000) | (tmp5999 & tmp6001) | (tmp6000 & tmp6001);
  wire tmp6003;
  assign tmp6003 = (tmp5994 & tmp5998) | (tmp5994 & tmp6002) | (tmp5998 & tmp6002);
  wire tmp6004;
  assign tmp6004 = 1'b1;
  wire tmp6005;
  assign tmp6005 = ~pi5;
  wire tmp6006;
  assign tmp6006 = ~pi6;
  wire tmp6007;
  assign tmp6007 = (tmp6004 & tmp6005) | (tmp6004 & tmp6006) | (tmp6005 & tmp6006);
  wire tmp6008;
  assign tmp6008 = ~pi5;
  wire tmp6009;
  assign tmp6009 = 1'b1;
  wire tmp6010;
  assign tmp6010 = 1'b1;
  wire tmp6011;
  assign tmp6011 = (tmp6008 & tmp6009) | (tmp6008 & tmp6010) | (tmp6009 & tmp6010);
  wire tmp6012;
  assign tmp6012 = ~pi6;
  wire tmp6013;
  assign tmp6013 = 1'b1;
  wire tmp6014;
  assign tmp6014 = 1'b1;
  wire tmp6015;
  assign tmp6015 = (tmp6012 & tmp6013) | (tmp6012 & tmp6014) | (tmp6013 & tmp6014);
  wire tmp6016;
  assign tmp6016 = (tmp6007 & tmp6011) | (tmp6007 & tmp6015) | (tmp6011 & tmp6015);
  wire tmp6017;
  assign tmp6017 = 1'b1;
  wire tmp6018;
  assign tmp6018 = ~pi6;
  wire tmp6019;
  assign tmp6019 = ~pi7;
  wire tmp6020;
  assign tmp6020 = (tmp6017 & tmp6018) | (tmp6017 & tmp6019) | (tmp6018 & tmp6019);
  wire tmp6021;
  assign tmp6021 = ~pi6;
  wire tmp6022;
  assign tmp6022 = 1'b1;
  wire tmp6023;
  assign tmp6023 = 1'b1;
  wire tmp6024;
  assign tmp6024 = (tmp6021 & tmp6022) | (tmp6021 & tmp6023) | (tmp6022 & tmp6023);
  wire tmp6025;
  assign tmp6025 = ~pi7;
  wire tmp6026;
  assign tmp6026 = 1'b1;
  wire tmp6027;
  assign tmp6027 = 1'b0;
  wire tmp6028;
  assign tmp6028 = (tmp6025 & tmp6026) | (tmp6025 & tmp6027) | (tmp6026 & tmp6027);
  wire tmp6029;
  assign tmp6029 = (tmp6020 & tmp6024) | (tmp6020 & tmp6028) | (tmp6024 & tmp6028);
  wire tmp6030;
  assign tmp6030 = (tmp6003 & tmp6016) | (tmp6003 & tmp6029) | (tmp6016 & tmp6029);
  wire tmp6031;
  assign tmp6031 = 1'b0;
  wire tmp6032;
  assign tmp6032 = 1'b1;
  wire tmp6033;
  assign tmp6033 = 1'b0;
  wire tmp6034;
  assign tmp6034 = (tmp6031 & tmp6032) | (tmp6031 & tmp6033) | (tmp6032 & tmp6033);
  wire tmp6035;
  assign tmp6035 = 1'b1;
  wire tmp6036;
  assign tmp6036 = ~pi6;
  wire tmp6037;
  assign tmp6037 = ~pi7;
  wire tmp6038;
  assign tmp6038 = (tmp6035 & tmp6036) | (tmp6035 & tmp6037) | (tmp6036 & tmp6037);
  wire tmp6039;
  assign tmp6039 = 1'b0;
  wire tmp6040;
  assign tmp6040 = ~pi7;
  wire tmp6041;
  assign tmp6041 = 1'b0;
  wire tmp6042;
  assign tmp6042 = (tmp6039 & tmp6040) | (tmp6039 & tmp6041) | (tmp6040 & tmp6041);
  wire tmp6043;
  assign tmp6043 = (tmp6034 & tmp6038) | (tmp6034 & tmp6042) | (tmp6038 & tmp6042);
  wire tmp6044;
  assign tmp6044 = 1'b1;
  wire tmp6045;
  assign tmp6045 = ~pi6;
  wire tmp6046;
  assign tmp6046 = ~pi7;
  wire tmp6047;
  assign tmp6047 = (tmp6044 & tmp6045) | (tmp6044 & tmp6046) | (tmp6045 & tmp6046);
  wire tmp6048;
  assign tmp6048 = ~pi6;
  wire tmp6049;
  assign tmp6049 = 1'b1;
  wire tmp6050;
  assign tmp6050 = 1'b1;
  wire tmp6051;
  assign tmp6051 = (tmp6048 & tmp6049) | (tmp6048 & tmp6050) | (tmp6049 & tmp6050);
  wire tmp6052;
  assign tmp6052 = ~pi7;
  wire tmp6053;
  assign tmp6053 = 1'b1;
  wire tmp6054;
  assign tmp6054 = 1'b0;
  wire tmp6055;
  assign tmp6055 = (tmp6052 & tmp6053) | (tmp6052 & tmp6054) | (tmp6053 & tmp6054);
  wire tmp6056;
  assign tmp6056 = (tmp6047 & tmp6051) | (tmp6047 & tmp6055) | (tmp6051 & tmp6055);
  wire tmp6057;
  assign tmp6057 = 1'b0;
  wire tmp6058;
  assign tmp6058 = ~pi7;
  wire tmp6059;
  assign tmp6059 = 1'b0;
  wire tmp6060;
  assign tmp6060 = (tmp6057 & tmp6058) | (tmp6057 & tmp6059) | (tmp6058 & tmp6059);
  wire tmp6061;
  assign tmp6061 = ~pi7;
  wire tmp6062;
  assign tmp6062 = 1'b1;
  wire tmp6063;
  assign tmp6063 = 1'b0;
  wire tmp6064;
  assign tmp6064 = (tmp6061 & tmp6062) | (tmp6061 & tmp6063) | (tmp6062 & tmp6063);
  wire tmp6065;
  assign tmp6065 = 1'b0;
  wire tmp6066;
  assign tmp6066 = 1'b0;
  wire tmp6067;
  assign tmp6067 = 1'b0;
  wire tmp6068;
  assign tmp6068 = (tmp6065 & tmp6066) | (tmp6065 & tmp6067) | (tmp6066 & tmp6067);
  wire tmp6069;
  assign tmp6069 = (tmp6060 & tmp6064) | (tmp6060 & tmp6068) | (tmp6064 & tmp6068);
  wire tmp6070;
  assign tmp6070 = (tmp6043 & tmp6056) | (tmp6043 & tmp6069) | (tmp6056 & tmp6069);
  wire tmp6071;
  assign tmp6071 = (tmp5990 & tmp6030) | (tmp5990 & tmp6070) | (tmp6030 & tmp6070);
  wire tmp6072;
  assign tmp6072 = 1'b0;
  wire tmp6073;
  assign tmp6073 = 1'b0;
  wire tmp6074;
  assign tmp6074 = 1'b0;
  wire tmp6075;
  assign tmp6075 = (tmp6072 & tmp6073) | (tmp6072 & tmp6074) | (tmp6073 & tmp6074);
  wire tmp6076;
  assign tmp6076 = 1'b0;
  wire tmp6077;
  assign tmp6077 = 1'b1;
  wire tmp6078;
  assign tmp6078 = 1'b0;
  wire tmp6079;
  assign tmp6079 = (tmp6076 & tmp6077) | (tmp6076 & tmp6078) | (tmp6077 & tmp6078);
  wire tmp6080;
  assign tmp6080 = 1'b0;
  wire tmp6081;
  assign tmp6081 = 1'b0;
  wire tmp6082;
  assign tmp6082 = 1'b0;
  wire tmp6083;
  assign tmp6083 = (tmp6080 & tmp6081) | (tmp6080 & tmp6082) | (tmp6081 & tmp6082);
  wire tmp6084;
  assign tmp6084 = (tmp6075 & tmp6079) | (tmp6075 & tmp6083) | (tmp6079 & tmp6083);
  wire tmp6085;
  assign tmp6085 = 1'b0;
  wire tmp6086;
  assign tmp6086 = 1'b1;
  wire tmp6087;
  assign tmp6087 = 1'b0;
  wire tmp6088;
  assign tmp6088 = (tmp6085 & tmp6086) | (tmp6085 & tmp6087) | (tmp6086 & tmp6087);
  wire tmp6089;
  assign tmp6089 = 1'b1;
  wire tmp6090;
  assign tmp6090 = ~pi6;
  wire tmp6091;
  assign tmp6091 = ~pi7;
  wire tmp6092;
  assign tmp6092 = (tmp6089 & tmp6090) | (tmp6089 & tmp6091) | (tmp6090 & tmp6091);
  wire tmp6093;
  assign tmp6093 = 1'b0;
  wire tmp6094;
  assign tmp6094 = ~pi7;
  wire tmp6095;
  assign tmp6095 = 1'b0;
  wire tmp6096;
  assign tmp6096 = (tmp6093 & tmp6094) | (tmp6093 & tmp6095) | (tmp6094 & tmp6095);
  wire tmp6097;
  assign tmp6097 = (tmp6088 & tmp6092) | (tmp6088 & tmp6096) | (tmp6092 & tmp6096);
  wire tmp6098;
  assign tmp6098 = 1'b0;
  wire tmp6099;
  assign tmp6099 = 1'b0;
  wire tmp6100;
  assign tmp6100 = 1'b0;
  wire tmp6101;
  assign tmp6101 = (tmp6098 & tmp6099) | (tmp6098 & tmp6100) | (tmp6099 & tmp6100);
  wire tmp6102;
  assign tmp6102 = 1'b0;
  wire tmp6103;
  assign tmp6103 = ~pi7;
  wire tmp6104;
  assign tmp6104 = 1'b0;
  wire tmp6105;
  assign tmp6105 = (tmp6102 & tmp6103) | (tmp6102 & tmp6104) | (tmp6103 & tmp6104);
  wire tmp6106;
  assign tmp6106 = 1'b0;
  wire tmp6107;
  assign tmp6107 = 1'b0;
  wire tmp6108;
  assign tmp6108 = 1'b0;
  wire tmp6109;
  assign tmp6109 = (tmp6106 & tmp6107) | (tmp6106 & tmp6108) | (tmp6107 & tmp6108);
  wire tmp6110;
  assign tmp6110 = (tmp6101 & tmp6105) | (tmp6101 & tmp6109) | (tmp6105 & tmp6109);
  wire tmp6111;
  assign tmp6111 = (tmp6084 & tmp6097) | (tmp6084 & tmp6110) | (tmp6097 & tmp6110);
  wire tmp6112;
  assign tmp6112 = 1'b0;
  wire tmp6113;
  assign tmp6113 = 1'b1;
  wire tmp6114;
  assign tmp6114 = 1'b0;
  wire tmp6115;
  assign tmp6115 = (tmp6112 & tmp6113) | (tmp6112 & tmp6114) | (tmp6113 & tmp6114);
  wire tmp6116;
  assign tmp6116 = 1'b1;
  wire tmp6117;
  assign tmp6117 = ~pi6;
  wire tmp6118;
  assign tmp6118 = ~pi7;
  wire tmp6119;
  assign tmp6119 = (tmp6116 & tmp6117) | (tmp6116 & tmp6118) | (tmp6117 & tmp6118);
  wire tmp6120;
  assign tmp6120 = 1'b0;
  wire tmp6121;
  assign tmp6121 = ~pi7;
  wire tmp6122;
  assign tmp6122 = 1'b0;
  wire tmp6123;
  assign tmp6123 = (tmp6120 & tmp6121) | (tmp6120 & tmp6122) | (tmp6121 & tmp6122);
  wire tmp6124;
  assign tmp6124 = (tmp6115 & tmp6119) | (tmp6115 & tmp6123) | (tmp6119 & tmp6123);
  wire tmp6125;
  assign tmp6125 = 1'b1;
  wire tmp6126;
  assign tmp6126 = ~pi6;
  wire tmp6127;
  assign tmp6127 = ~pi7;
  wire tmp6128;
  assign tmp6128 = (tmp6125 & tmp6126) | (tmp6125 & tmp6127) | (tmp6126 & tmp6127);
  wire tmp6129;
  assign tmp6129 = ~pi6;
  wire tmp6130;
  assign tmp6130 = 1'b1;
  wire tmp6131;
  assign tmp6131 = 1'b1;
  wire tmp6132;
  assign tmp6132 = (tmp6129 & tmp6130) | (tmp6129 & tmp6131) | (tmp6130 & tmp6131);
  wire tmp6133;
  assign tmp6133 = ~pi7;
  wire tmp6134;
  assign tmp6134 = 1'b1;
  wire tmp6135;
  assign tmp6135 = 1'b0;
  wire tmp6136;
  assign tmp6136 = (tmp6133 & tmp6134) | (tmp6133 & tmp6135) | (tmp6134 & tmp6135);
  wire tmp6137;
  assign tmp6137 = (tmp6128 & tmp6132) | (tmp6128 & tmp6136) | (tmp6132 & tmp6136);
  wire tmp6138;
  assign tmp6138 = 1'b0;
  wire tmp6139;
  assign tmp6139 = ~pi7;
  wire tmp6140;
  assign tmp6140 = 1'b0;
  wire tmp6141;
  assign tmp6141 = (tmp6138 & tmp6139) | (tmp6138 & tmp6140) | (tmp6139 & tmp6140);
  wire tmp6142;
  assign tmp6142 = ~pi7;
  wire tmp6143;
  assign tmp6143 = 1'b1;
  wire tmp6144;
  assign tmp6144 = 1'b0;
  wire tmp6145;
  assign tmp6145 = (tmp6142 & tmp6143) | (tmp6142 & tmp6144) | (tmp6143 & tmp6144);
  wire tmp6146;
  assign tmp6146 = 1'b0;
  wire tmp6147;
  assign tmp6147 = 1'b0;
  wire tmp6148;
  assign tmp6148 = 1'b0;
  wire tmp6149;
  assign tmp6149 = (tmp6146 & tmp6147) | (tmp6146 & tmp6148) | (tmp6147 & tmp6148);
  wire tmp6150;
  assign tmp6150 = (tmp6141 & tmp6145) | (tmp6141 & tmp6149) | (tmp6145 & tmp6149);
  wire tmp6151;
  assign tmp6151 = (tmp6124 & tmp6137) | (tmp6124 & tmp6150) | (tmp6137 & tmp6150);
  wire tmp6152;
  assign tmp6152 = 1'b0;
  wire tmp6153;
  assign tmp6153 = 1'b0;
  wire tmp6154;
  assign tmp6154 = 1'b0;
  wire tmp6155;
  assign tmp6155 = (tmp6152 & tmp6153) | (tmp6152 & tmp6154) | (tmp6153 & tmp6154);
  wire tmp6156;
  assign tmp6156 = 1'b0;
  wire tmp6157;
  assign tmp6157 = ~pi7;
  wire tmp6158;
  assign tmp6158 = 1'b0;
  wire tmp6159;
  assign tmp6159 = (tmp6156 & tmp6157) | (tmp6156 & tmp6158) | (tmp6157 & tmp6158);
  wire tmp6160;
  assign tmp6160 = 1'b0;
  wire tmp6161;
  assign tmp6161 = 1'b0;
  wire tmp6162;
  assign tmp6162 = 1'b0;
  wire tmp6163;
  assign tmp6163 = (tmp6160 & tmp6161) | (tmp6160 & tmp6162) | (tmp6161 & tmp6162);
  wire tmp6164;
  assign tmp6164 = (tmp6155 & tmp6159) | (tmp6155 & tmp6163) | (tmp6159 & tmp6163);
  wire tmp6165;
  assign tmp6165 = 1'b0;
  wire tmp6166;
  assign tmp6166 = ~pi7;
  wire tmp6167;
  assign tmp6167 = 1'b0;
  wire tmp6168;
  assign tmp6168 = (tmp6165 & tmp6166) | (tmp6165 & tmp6167) | (tmp6166 & tmp6167);
  wire tmp6169;
  assign tmp6169 = ~pi7;
  wire tmp6170;
  assign tmp6170 = 1'b1;
  wire tmp6171;
  assign tmp6171 = 1'b0;
  wire tmp6172;
  assign tmp6172 = (tmp6169 & tmp6170) | (tmp6169 & tmp6171) | (tmp6170 & tmp6171);
  wire tmp6173;
  assign tmp6173 = 1'b0;
  wire tmp6174;
  assign tmp6174 = 1'b0;
  wire tmp6175;
  assign tmp6175 = 1'b0;
  wire tmp6176;
  assign tmp6176 = (tmp6173 & tmp6174) | (tmp6173 & tmp6175) | (tmp6174 & tmp6175);
  wire tmp6177;
  assign tmp6177 = (tmp6168 & tmp6172) | (tmp6168 & tmp6176) | (tmp6172 & tmp6176);
  wire tmp6178;
  assign tmp6178 = 1'b0;
  wire tmp6179;
  assign tmp6179 = 1'b0;
  wire tmp6180;
  assign tmp6180 = 1'b0;
  wire tmp6181;
  assign tmp6181 = (tmp6178 & tmp6179) | (tmp6178 & tmp6180) | (tmp6179 & tmp6180);
  wire tmp6182;
  assign tmp6182 = 1'b0;
  wire tmp6183;
  assign tmp6183 = 1'b0;
  wire tmp6184;
  assign tmp6184 = 1'b0;
  wire tmp6185;
  assign tmp6185 = (tmp6182 & tmp6183) | (tmp6182 & tmp6184) | (tmp6183 & tmp6184);
  wire tmp6186;
  assign tmp6186 = 1'b0;
  wire tmp6187;
  assign tmp6187 = 1'b0;
  wire tmp6188;
  assign tmp6188 = 1'b0;
  wire tmp6189;
  assign tmp6189 = (tmp6186 & tmp6187) | (tmp6186 & tmp6188) | (tmp6187 & tmp6188);
  wire tmp6190;
  assign tmp6190 = (tmp6181 & tmp6185) | (tmp6181 & tmp6189) | (tmp6185 & tmp6189);
  wire tmp6191;
  assign tmp6191 = (tmp6164 & tmp6177) | (tmp6164 & tmp6190) | (tmp6177 & tmp6190);
  wire tmp6192;
  assign tmp6192 = (tmp6111 & tmp6151) | (tmp6111 & tmp6191) | (tmp6151 & tmp6191);
  wire tmp6193;
  assign tmp6193 = (tmp5950 & tmp6071) | (tmp5950 & tmp6192) | (tmp6071 & tmp6192);
  wire tmp6194;
  assign tmp6194 = 1'b0;
  wire tmp6195;
  assign tmp6195 = 1'b0;
  wire tmp6196;
  assign tmp6196 = 1'b0;
  wire tmp6197;
  assign tmp6197 = (tmp6194 & tmp6195) | (tmp6194 & tmp6196) | (tmp6195 & tmp6196);
  wire tmp6198;
  assign tmp6198 = 1'b0;
  wire tmp6199;
  assign tmp6199 = 1'b0;
  wire tmp6200;
  assign tmp6200 = 1'b0;
  wire tmp6201;
  assign tmp6201 = (tmp6198 & tmp6199) | (tmp6198 & tmp6200) | (tmp6199 & tmp6200);
  wire tmp6202;
  assign tmp6202 = 1'b0;
  wire tmp6203;
  assign tmp6203 = 1'b0;
  wire tmp6204;
  assign tmp6204 = 1'b0;
  wire tmp6205;
  assign tmp6205 = (tmp6202 & tmp6203) | (tmp6202 & tmp6204) | (tmp6203 & tmp6204);
  wire tmp6206;
  assign tmp6206 = (tmp6197 & tmp6201) | (tmp6197 & tmp6205) | (tmp6201 & tmp6205);
  wire tmp6207;
  assign tmp6207 = 1'b0;
  wire tmp6208;
  assign tmp6208 = 1'b0;
  wire tmp6209;
  assign tmp6209 = 1'b0;
  wire tmp6210;
  assign tmp6210 = (tmp6207 & tmp6208) | (tmp6207 & tmp6209) | (tmp6208 & tmp6209);
  wire tmp6211;
  assign tmp6211 = 1'b0;
  wire tmp6212;
  assign tmp6212 = 1'b1;
  wire tmp6213;
  assign tmp6213 = 1'b0;
  wire tmp6214;
  assign tmp6214 = (tmp6211 & tmp6212) | (tmp6211 & tmp6213) | (tmp6212 & tmp6213);
  wire tmp6215;
  assign tmp6215 = 1'b0;
  wire tmp6216;
  assign tmp6216 = 1'b0;
  wire tmp6217;
  assign tmp6217 = 1'b0;
  wire tmp6218;
  assign tmp6218 = (tmp6215 & tmp6216) | (tmp6215 & tmp6217) | (tmp6216 & tmp6217);
  wire tmp6219;
  assign tmp6219 = (tmp6210 & tmp6214) | (tmp6210 & tmp6218) | (tmp6214 & tmp6218);
  wire tmp6220;
  assign tmp6220 = 1'b0;
  wire tmp6221;
  assign tmp6221 = 1'b0;
  wire tmp6222;
  assign tmp6222 = 1'b0;
  wire tmp6223;
  assign tmp6223 = (tmp6220 & tmp6221) | (tmp6220 & tmp6222) | (tmp6221 & tmp6222);
  wire tmp6224;
  assign tmp6224 = 1'b0;
  wire tmp6225;
  assign tmp6225 = 1'b0;
  wire tmp6226;
  assign tmp6226 = 1'b0;
  wire tmp6227;
  assign tmp6227 = (tmp6224 & tmp6225) | (tmp6224 & tmp6226) | (tmp6225 & tmp6226);
  wire tmp6228;
  assign tmp6228 = 1'b0;
  wire tmp6229;
  assign tmp6229 = 1'b0;
  wire tmp6230;
  assign tmp6230 = 1'b0;
  wire tmp6231;
  assign tmp6231 = (tmp6228 & tmp6229) | (tmp6228 & tmp6230) | (tmp6229 & tmp6230);
  wire tmp6232;
  assign tmp6232 = (tmp6223 & tmp6227) | (tmp6223 & tmp6231) | (tmp6227 & tmp6231);
  wire tmp6233;
  assign tmp6233 = (tmp6206 & tmp6219) | (tmp6206 & tmp6232) | (tmp6219 & tmp6232);
  wire tmp6234;
  assign tmp6234 = 1'b0;
  wire tmp6235;
  assign tmp6235 = 1'b0;
  wire tmp6236;
  assign tmp6236 = 1'b0;
  wire tmp6237;
  assign tmp6237 = (tmp6234 & tmp6235) | (tmp6234 & tmp6236) | (tmp6235 & tmp6236);
  wire tmp6238;
  assign tmp6238 = 1'b0;
  wire tmp6239;
  assign tmp6239 = 1'b1;
  wire tmp6240;
  assign tmp6240 = 1'b0;
  wire tmp6241;
  assign tmp6241 = (tmp6238 & tmp6239) | (tmp6238 & tmp6240) | (tmp6239 & tmp6240);
  wire tmp6242;
  assign tmp6242 = 1'b0;
  wire tmp6243;
  assign tmp6243 = 1'b0;
  wire tmp6244;
  assign tmp6244 = 1'b0;
  wire tmp6245;
  assign tmp6245 = (tmp6242 & tmp6243) | (tmp6242 & tmp6244) | (tmp6243 & tmp6244);
  wire tmp6246;
  assign tmp6246 = (tmp6237 & tmp6241) | (tmp6237 & tmp6245) | (tmp6241 & tmp6245);
  wire tmp6247;
  assign tmp6247 = 1'b0;
  wire tmp6248;
  assign tmp6248 = 1'b1;
  wire tmp6249;
  assign tmp6249 = 1'b0;
  wire tmp6250;
  assign tmp6250 = (tmp6247 & tmp6248) | (tmp6247 & tmp6249) | (tmp6248 & tmp6249);
  wire tmp6251;
  assign tmp6251 = 1'b1;
  wire tmp6252;
  assign tmp6252 = ~pi6;
  wire tmp6253;
  assign tmp6253 = ~pi7;
  wire tmp6254;
  assign tmp6254 = (tmp6251 & tmp6252) | (tmp6251 & tmp6253) | (tmp6252 & tmp6253);
  wire tmp6255;
  assign tmp6255 = 1'b0;
  wire tmp6256;
  assign tmp6256 = ~pi7;
  wire tmp6257;
  assign tmp6257 = 1'b0;
  wire tmp6258;
  assign tmp6258 = (tmp6255 & tmp6256) | (tmp6255 & tmp6257) | (tmp6256 & tmp6257);
  wire tmp6259;
  assign tmp6259 = (tmp6250 & tmp6254) | (tmp6250 & tmp6258) | (tmp6254 & tmp6258);
  wire tmp6260;
  assign tmp6260 = 1'b0;
  wire tmp6261;
  assign tmp6261 = 1'b0;
  wire tmp6262;
  assign tmp6262 = 1'b0;
  wire tmp6263;
  assign tmp6263 = (tmp6260 & tmp6261) | (tmp6260 & tmp6262) | (tmp6261 & tmp6262);
  wire tmp6264;
  assign tmp6264 = 1'b0;
  wire tmp6265;
  assign tmp6265 = ~pi7;
  wire tmp6266;
  assign tmp6266 = 1'b0;
  wire tmp6267;
  assign tmp6267 = (tmp6264 & tmp6265) | (tmp6264 & tmp6266) | (tmp6265 & tmp6266);
  wire tmp6268;
  assign tmp6268 = 1'b0;
  wire tmp6269;
  assign tmp6269 = 1'b0;
  wire tmp6270;
  assign tmp6270 = 1'b0;
  wire tmp6271;
  assign tmp6271 = (tmp6268 & tmp6269) | (tmp6268 & tmp6270) | (tmp6269 & tmp6270);
  wire tmp6272;
  assign tmp6272 = (tmp6263 & tmp6267) | (tmp6263 & tmp6271) | (tmp6267 & tmp6271);
  wire tmp6273;
  assign tmp6273 = (tmp6246 & tmp6259) | (tmp6246 & tmp6272) | (tmp6259 & tmp6272);
  wire tmp6274;
  assign tmp6274 = 1'b0;
  wire tmp6275;
  assign tmp6275 = 1'b0;
  wire tmp6276;
  assign tmp6276 = 1'b0;
  wire tmp6277;
  assign tmp6277 = (tmp6274 & tmp6275) | (tmp6274 & tmp6276) | (tmp6275 & tmp6276);
  wire tmp6278;
  assign tmp6278 = 1'b0;
  wire tmp6279;
  assign tmp6279 = 1'b0;
  wire tmp6280;
  assign tmp6280 = 1'b0;
  wire tmp6281;
  assign tmp6281 = (tmp6278 & tmp6279) | (tmp6278 & tmp6280) | (tmp6279 & tmp6280);
  wire tmp6282;
  assign tmp6282 = 1'b0;
  wire tmp6283;
  assign tmp6283 = 1'b0;
  wire tmp6284;
  assign tmp6284 = 1'b0;
  wire tmp6285;
  assign tmp6285 = (tmp6282 & tmp6283) | (tmp6282 & tmp6284) | (tmp6283 & tmp6284);
  wire tmp6286;
  assign tmp6286 = (tmp6277 & tmp6281) | (tmp6277 & tmp6285) | (tmp6281 & tmp6285);
  wire tmp6287;
  assign tmp6287 = 1'b0;
  wire tmp6288;
  assign tmp6288 = 1'b0;
  wire tmp6289;
  assign tmp6289 = 1'b0;
  wire tmp6290;
  assign tmp6290 = (tmp6287 & tmp6288) | (tmp6287 & tmp6289) | (tmp6288 & tmp6289);
  wire tmp6291;
  assign tmp6291 = 1'b0;
  wire tmp6292;
  assign tmp6292 = ~pi7;
  wire tmp6293;
  assign tmp6293 = 1'b0;
  wire tmp6294;
  assign tmp6294 = (tmp6291 & tmp6292) | (tmp6291 & tmp6293) | (tmp6292 & tmp6293);
  wire tmp6295;
  assign tmp6295 = 1'b0;
  wire tmp6296;
  assign tmp6296 = 1'b0;
  wire tmp6297;
  assign tmp6297 = 1'b0;
  wire tmp6298;
  assign tmp6298 = (tmp6295 & tmp6296) | (tmp6295 & tmp6297) | (tmp6296 & tmp6297);
  wire tmp6299;
  assign tmp6299 = (tmp6290 & tmp6294) | (tmp6290 & tmp6298) | (tmp6294 & tmp6298);
  wire tmp6300;
  assign tmp6300 = 1'b0;
  wire tmp6301;
  assign tmp6301 = 1'b0;
  wire tmp6302;
  assign tmp6302 = 1'b0;
  wire tmp6303;
  assign tmp6303 = (tmp6300 & tmp6301) | (tmp6300 & tmp6302) | (tmp6301 & tmp6302);
  wire tmp6304;
  assign tmp6304 = 1'b0;
  wire tmp6305;
  assign tmp6305 = 1'b0;
  wire tmp6306;
  assign tmp6306 = 1'b0;
  wire tmp6307;
  assign tmp6307 = (tmp6304 & tmp6305) | (tmp6304 & tmp6306) | (tmp6305 & tmp6306);
  wire tmp6308;
  assign tmp6308 = 1'b0;
  wire tmp6309;
  assign tmp6309 = 1'b0;
  wire tmp6310;
  assign tmp6310 = 1'b0;
  wire tmp6311;
  assign tmp6311 = (tmp6308 & tmp6309) | (tmp6308 & tmp6310) | (tmp6309 & tmp6310);
  wire tmp6312;
  assign tmp6312 = (tmp6303 & tmp6307) | (tmp6303 & tmp6311) | (tmp6307 & tmp6311);
  wire tmp6313;
  assign tmp6313 = (tmp6286 & tmp6299) | (tmp6286 & tmp6312) | (tmp6299 & tmp6312);
  wire tmp6314;
  assign tmp6314 = (tmp6233 & tmp6273) | (tmp6233 & tmp6313) | (tmp6273 & tmp6313);
  wire tmp6315;
  assign tmp6315 = 1'b0;
  wire tmp6316;
  assign tmp6316 = 1'b0;
  wire tmp6317;
  assign tmp6317 = 1'b0;
  wire tmp6318;
  assign tmp6318 = (tmp6315 & tmp6316) | (tmp6315 & tmp6317) | (tmp6316 & tmp6317);
  wire tmp6319;
  assign tmp6319 = 1'b0;
  wire tmp6320;
  assign tmp6320 = 1'b1;
  wire tmp6321;
  assign tmp6321 = 1'b0;
  wire tmp6322;
  assign tmp6322 = (tmp6319 & tmp6320) | (tmp6319 & tmp6321) | (tmp6320 & tmp6321);
  wire tmp6323;
  assign tmp6323 = 1'b0;
  wire tmp6324;
  assign tmp6324 = 1'b0;
  wire tmp6325;
  assign tmp6325 = 1'b0;
  wire tmp6326;
  assign tmp6326 = (tmp6323 & tmp6324) | (tmp6323 & tmp6325) | (tmp6324 & tmp6325);
  wire tmp6327;
  assign tmp6327 = (tmp6318 & tmp6322) | (tmp6318 & tmp6326) | (tmp6322 & tmp6326);
  wire tmp6328;
  assign tmp6328 = 1'b0;
  wire tmp6329;
  assign tmp6329 = 1'b1;
  wire tmp6330;
  assign tmp6330 = 1'b0;
  wire tmp6331;
  assign tmp6331 = (tmp6328 & tmp6329) | (tmp6328 & tmp6330) | (tmp6329 & tmp6330);
  wire tmp6332;
  assign tmp6332 = 1'b1;
  wire tmp6333;
  assign tmp6333 = ~pi6;
  wire tmp6334;
  assign tmp6334 = ~pi7;
  wire tmp6335;
  assign tmp6335 = (tmp6332 & tmp6333) | (tmp6332 & tmp6334) | (tmp6333 & tmp6334);
  wire tmp6336;
  assign tmp6336 = 1'b0;
  wire tmp6337;
  assign tmp6337 = ~pi7;
  wire tmp6338;
  assign tmp6338 = 1'b0;
  wire tmp6339;
  assign tmp6339 = (tmp6336 & tmp6337) | (tmp6336 & tmp6338) | (tmp6337 & tmp6338);
  wire tmp6340;
  assign tmp6340 = (tmp6331 & tmp6335) | (tmp6331 & tmp6339) | (tmp6335 & tmp6339);
  wire tmp6341;
  assign tmp6341 = 1'b0;
  wire tmp6342;
  assign tmp6342 = 1'b0;
  wire tmp6343;
  assign tmp6343 = 1'b0;
  wire tmp6344;
  assign tmp6344 = (tmp6341 & tmp6342) | (tmp6341 & tmp6343) | (tmp6342 & tmp6343);
  wire tmp6345;
  assign tmp6345 = 1'b0;
  wire tmp6346;
  assign tmp6346 = ~pi7;
  wire tmp6347;
  assign tmp6347 = 1'b0;
  wire tmp6348;
  assign tmp6348 = (tmp6345 & tmp6346) | (tmp6345 & tmp6347) | (tmp6346 & tmp6347);
  wire tmp6349;
  assign tmp6349 = 1'b0;
  wire tmp6350;
  assign tmp6350 = 1'b0;
  wire tmp6351;
  assign tmp6351 = 1'b0;
  wire tmp6352;
  assign tmp6352 = (tmp6349 & tmp6350) | (tmp6349 & tmp6351) | (tmp6350 & tmp6351);
  wire tmp6353;
  assign tmp6353 = (tmp6344 & tmp6348) | (tmp6344 & tmp6352) | (tmp6348 & tmp6352);
  wire tmp6354;
  assign tmp6354 = (tmp6327 & tmp6340) | (tmp6327 & tmp6353) | (tmp6340 & tmp6353);
  wire tmp6355;
  assign tmp6355 = 1'b0;
  wire tmp6356;
  assign tmp6356 = 1'b1;
  wire tmp6357;
  assign tmp6357 = 1'b0;
  wire tmp6358;
  assign tmp6358 = (tmp6355 & tmp6356) | (tmp6355 & tmp6357) | (tmp6356 & tmp6357);
  wire tmp6359;
  assign tmp6359 = 1'b1;
  wire tmp6360;
  assign tmp6360 = ~pi6;
  wire tmp6361;
  assign tmp6361 = ~pi7;
  wire tmp6362;
  assign tmp6362 = (tmp6359 & tmp6360) | (tmp6359 & tmp6361) | (tmp6360 & tmp6361);
  wire tmp6363;
  assign tmp6363 = 1'b0;
  wire tmp6364;
  assign tmp6364 = ~pi7;
  wire tmp6365;
  assign tmp6365 = 1'b0;
  wire tmp6366;
  assign tmp6366 = (tmp6363 & tmp6364) | (tmp6363 & tmp6365) | (tmp6364 & tmp6365);
  wire tmp6367;
  assign tmp6367 = (tmp6358 & tmp6362) | (tmp6358 & tmp6366) | (tmp6362 & tmp6366);
  wire tmp6368;
  assign tmp6368 = 1'b1;
  wire tmp6369;
  assign tmp6369 = ~pi6;
  wire tmp6370;
  assign tmp6370 = ~pi7;
  wire tmp6371;
  assign tmp6371 = (tmp6368 & tmp6369) | (tmp6368 & tmp6370) | (tmp6369 & tmp6370);
  wire tmp6372;
  assign tmp6372 = ~pi6;
  wire tmp6373;
  assign tmp6373 = 1'b1;
  wire tmp6374;
  assign tmp6374 = 1'b1;
  wire tmp6375;
  assign tmp6375 = (tmp6372 & tmp6373) | (tmp6372 & tmp6374) | (tmp6373 & tmp6374);
  wire tmp6376;
  assign tmp6376 = ~pi7;
  wire tmp6377;
  assign tmp6377 = 1'b1;
  wire tmp6378;
  assign tmp6378 = 1'b0;
  wire tmp6379;
  assign tmp6379 = (tmp6376 & tmp6377) | (tmp6376 & tmp6378) | (tmp6377 & tmp6378);
  wire tmp6380;
  assign tmp6380 = (tmp6371 & tmp6375) | (tmp6371 & tmp6379) | (tmp6375 & tmp6379);
  wire tmp6381;
  assign tmp6381 = 1'b0;
  wire tmp6382;
  assign tmp6382 = ~pi7;
  wire tmp6383;
  assign tmp6383 = 1'b0;
  wire tmp6384;
  assign tmp6384 = (tmp6381 & tmp6382) | (tmp6381 & tmp6383) | (tmp6382 & tmp6383);
  wire tmp6385;
  assign tmp6385 = ~pi7;
  wire tmp6386;
  assign tmp6386 = 1'b1;
  wire tmp6387;
  assign tmp6387 = 1'b0;
  wire tmp6388;
  assign tmp6388 = (tmp6385 & tmp6386) | (tmp6385 & tmp6387) | (tmp6386 & tmp6387);
  wire tmp6389;
  assign tmp6389 = 1'b0;
  wire tmp6390;
  assign tmp6390 = 1'b0;
  wire tmp6391;
  assign tmp6391 = 1'b0;
  wire tmp6392;
  assign tmp6392 = (tmp6389 & tmp6390) | (tmp6389 & tmp6391) | (tmp6390 & tmp6391);
  wire tmp6393;
  assign tmp6393 = (tmp6384 & tmp6388) | (tmp6384 & tmp6392) | (tmp6388 & tmp6392);
  wire tmp6394;
  assign tmp6394 = (tmp6367 & tmp6380) | (tmp6367 & tmp6393) | (tmp6380 & tmp6393);
  wire tmp6395;
  assign tmp6395 = 1'b0;
  wire tmp6396;
  assign tmp6396 = 1'b0;
  wire tmp6397;
  assign tmp6397 = 1'b0;
  wire tmp6398;
  assign tmp6398 = (tmp6395 & tmp6396) | (tmp6395 & tmp6397) | (tmp6396 & tmp6397);
  wire tmp6399;
  assign tmp6399 = 1'b0;
  wire tmp6400;
  assign tmp6400 = ~pi7;
  wire tmp6401;
  assign tmp6401 = 1'b0;
  wire tmp6402;
  assign tmp6402 = (tmp6399 & tmp6400) | (tmp6399 & tmp6401) | (tmp6400 & tmp6401);
  wire tmp6403;
  assign tmp6403 = 1'b0;
  wire tmp6404;
  assign tmp6404 = 1'b0;
  wire tmp6405;
  assign tmp6405 = 1'b0;
  wire tmp6406;
  assign tmp6406 = (tmp6403 & tmp6404) | (tmp6403 & tmp6405) | (tmp6404 & tmp6405);
  wire tmp6407;
  assign tmp6407 = (tmp6398 & tmp6402) | (tmp6398 & tmp6406) | (tmp6402 & tmp6406);
  wire tmp6408;
  assign tmp6408 = 1'b0;
  wire tmp6409;
  assign tmp6409 = ~pi7;
  wire tmp6410;
  assign tmp6410 = 1'b0;
  wire tmp6411;
  assign tmp6411 = (tmp6408 & tmp6409) | (tmp6408 & tmp6410) | (tmp6409 & tmp6410);
  wire tmp6412;
  assign tmp6412 = ~pi7;
  wire tmp6413;
  assign tmp6413 = 1'b1;
  wire tmp6414;
  assign tmp6414 = 1'b0;
  wire tmp6415;
  assign tmp6415 = (tmp6412 & tmp6413) | (tmp6412 & tmp6414) | (tmp6413 & tmp6414);
  wire tmp6416;
  assign tmp6416 = 1'b0;
  wire tmp6417;
  assign tmp6417 = 1'b0;
  wire tmp6418;
  assign tmp6418 = 1'b0;
  wire tmp6419;
  assign tmp6419 = (tmp6416 & tmp6417) | (tmp6416 & tmp6418) | (tmp6417 & tmp6418);
  wire tmp6420;
  assign tmp6420 = (tmp6411 & tmp6415) | (tmp6411 & tmp6419) | (tmp6415 & tmp6419);
  wire tmp6421;
  assign tmp6421 = 1'b0;
  wire tmp6422;
  assign tmp6422 = 1'b0;
  wire tmp6423;
  assign tmp6423 = 1'b0;
  wire tmp6424;
  assign tmp6424 = (tmp6421 & tmp6422) | (tmp6421 & tmp6423) | (tmp6422 & tmp6423);
  wire tmp6425;
  assign tmp6425 = 1'b0;
  wire tmp6426;
  assign tmp6426 = 1'b0;
  wire tmp6427;
  assign tmp6427 = 1'b0;
  wire tmp6428;
  assign tmp6428 = (tmp6425 & tmp6426) | (tmp6425 & tmp6427) | (tmp6426 & tmp6427);
  wire tmp6429;
  assign tmp6429 = 1'b0;
  wire tmp6430;
  assign tmp6430 = 1'b0;
  wire tmp6431;
  assign tmp6431 = 1'b0;
  wire tmp6432;
  assign tmp6432 = (tmp6429 & tmp6430) | (tmp6429 & tmp6431) | (tmp6430 & tmp6431);
  wire tmp6433;
  assign tmp6433 = (tmp6424 & tmp6428) | (tmp6424 & tmp6432) | (tmp6428 & tmp6432);
  wire tmp6434;
  assign tmp6434 = (tmp6407 & tmp6420) | (tmp6407 & tmp6433) | (tmp6420 & tmp6433);
  wire tmp6435;
  assign tmp6435 = (tmp6354 & tmp6394) | (tmp6354 & tmp6434) | (tmp6394 & tmp6434);
  wire tmp6436;
  assign tmp6436 = 1'b0;
  wire tmp6437;
  assign tmp6437 = 1'b0;
  wire tmp6438;
  assign tmp6438 = 1'b0;
  wire tmp6439;
  assign tmp6439 = (tmp6436 & tmp6437) | (tmp6436 & tmp6438) | (tmp6437 & tmp6438);
  wire tmp6440;
  assign tmp6440 = 1'b0;
  wire tmp6441;
  assign tmp6441 = 1'b0;
  wire tmp6442;
  assign tmp6442 = 1'b0;
  wire tmp6443;
  assign tmp6443 = (tmp6440 & tmp6441) | (tmp6440 & tmp6442) | (tmp6441 & tmp6442);
  wire tmp6444;
  assign tmp6444 = 1'b0;
  wire tmp6445;
  assign tmp6445 = 1'b0;
  wire tmp6446;
  assign tmp6446 = 1'b0;
  wire tmp6447;
  assign tmp6447 = (tmp6444 & tmp6445) | (tmp6444 & tmp6446) | (tmp6445 & tmp6446);
  wire tmp6448;
  assign tmp6448 = (tmp6439 & tmp6443) | (tmp6439 & tmp6447) | (tmp6443 & tmp6447);
  wire tmp6449;
  assign tmp6449 = 1'b0;
  wire tmp6450;
  assign tmp6450 = 1'b0;
  wire tmp6451;
  assign tmp6451 = 1'b0;
  wire tmp6452;
  assign tmp6452 = (tmp6449 & tmp6450) | (tmp6449 & tmp6451) | (tmp6450 & tmp6451);
  wire tmp6453;
  assign tmp6453 = 1'b0;
  wire tmp6454;
  assign tmp6454 = ~pi7;
  wire tmp6455;
  assign tmp6455 = 1'b0;
  wire tmp6456;
  assign tmp6456 = (tmp6453 & tmp6454) | (tmp6453 & tmp6455) | (tmp6454 & tmp6455);
  wire tmp6457;
  assign tmp6457 = 1'b0;
  wire tmp6458;
  assign tmp6458 = 1'b0;
  wire tmp6459;
  assign tmp6459 = 1'b0;
  wire tmp6460;
  assign tmp6460 = (tmp6457 & tmp6458) | (tmp6457 & tmp6459) | (tmp6458 & tmp6459);
  wire tmp6461;
  assign tmp6461 = (tmp6452 & tmp6456) | (tmp6452 & tmp6460) | (tmp6456 & tmp6460);
  wire tmp6462;
  assign tmp6462 = 1'b0;
  wire tmp6463;
  assign tmp6463 = 1'b0;
  wire tmp6464;
  assign tmp6464 = 1'b0;
  wire tmp6465;
  assign tmp6465 = (tmp6462 & tmp6463) | (tmp6462 & tmp6464) | (tmp6463 & tmp6464);
  wire tmp6466;
  assign tmp6466 = 1'b0;
  wire tmp6467;
  assign tmp6467 = 1'b0;
  wire tmp6468;
  assign tmp6468 = 1'b0;
  wire tmp6469;
  assign tmp6469 = (tmp6466 & tmp6467) | (tmp6466 & tmp6468) | (tmp6467 & tmp6468);
  wire tmp6470;
  assign tmp6470 = 1'b0;
  wire tmp6471;
  assign tmp6471 = 1'b0;
  wire tmp6472;
  assign tmp6472 = 1'b0;
  wire tmp6473;
  assign tmp6473 = (tmp6470 & tmp6471) | (tmp6470 & tmp6472) | (tmp6471 & tmp6472);
  wire tmp6474;
  assign tmp6474 = (tmp6465 & tmp6469) | (tmp6465 & tmp6473) | (tmp6469 & tmp6473);
  wire tmp6475;
  assign tmp6475 = (tmp6448 & tmp6461) | (tmp6448 & tmp6474) | (tmp6461 & tmp6474);
  wire tmp6476;
  assign tmp6476 = 1'b0;
  wire tmp6477;
  assign tmp6477 = 1'b0;
  wire tmp6478;
  assign tmp6478 = 1'b0;
  wire tmp6479;
  assign tmp6479 = (tmp6476 & tmp6477) | (tmp6476 & tmp6478) | (tmp6477 & tmp6478);
  wire tmp6480;
  assign tmp6480 = 1'b0;
  wire tmp6481;
  assign tmp6481 = ~pi7;
  wire tmp6482;
  assign tmp6482 = 1'b0;
  wire tmp6483;
  assign tmp6483 = (tmp6480 & tmp6481) | (tmp6480 & tmp6482) | (tmp6481 & tmp6482);
  wire tmp6484;
  assign tmp6484 = 1'b0;
  wire tmp6485;
  assign tmp6485 = 1'b0;
  wire tmp6486;
  assign tmp6486 = 1'b0;
  wire tmp6487;
  assign tmp6487 = (tmp6484 & tmp6485) | (tmp6484 & tmp6486) | (tmp6485 & tmp6486);
  wire tmp6488;
  assign tmp6488 = (tmp6479 & tmp6483) | (tmp6479 & tmp6487) | (tmp6483 & tmp6487);
  wire tmp6489;
  assign tmp6489 = 1'b0;
  wire tmp6490;
  assign tmp6490 = ~pi7;
  wire tmp6491;
  assign tmp6491 = 1'b0;
  wire tmp6492;
  assign tmp6492 = (tmp6489 & tmp6490) | (tmp6489 & tmp6491) | (tmp6490 & tmp6491);
  wire tmp6493;
  assign tmp6493 = ~pi7;
  wire tmp6494;
  assign tmp6494 = 1'b1;
  wire tmp6495;
  assign tmp6495 = 1'b0;
  wire tmp6496;
  assign tmp6496 = (tmp6493 & tmp6494) | (tmp6493 & tmp6495) | (tmp6494 & tmp6495);
  wire tmp6497;
  assign tmp6497 = 1'b0;
  wire tmp6498;
  assign tmp6498 = 1'b0;
  wire tmp6499;
  assign tmp6499 = 1'b0;
  wire tmp6500;
  assign tmp6500 = (tmp6497 & tmp6498) | (tmp6497 & tmp6499) | (tmp6498 & tmp6499);
  wire tmp6501;
  assign tmp6501 = (tmp6492 & tmp6496) | (tmp6492 & tmp6500) | (tmp6496 & tmp6500);
  wire tmp6502;
  assign tmp6502 = 1'b0;
  wire tmp6503;
  assign tmp6503 = 1'b0;
  wire tmp6504;
  assign tmp6504 = 1'b0;
  wire tmp6505;
  assign tmp6505 = (tmp6502 & tmp6503) | (tmp6502 & tmp6504) | (tmp6503 & tmp6504);
  wire tmp6506;
  assign tmp6506 = 1'b0;
  wire tmp6507;
  assign tmp6507 = 1'b0;
  wire tmp6508;
  assign tmp6508 = 1'b0;
  wire tmp6509;
  assign tmp6509 = (tmp6506 & tmp6507) | (tmp6506 & tmp6508) | (tmp6507 & tmp6508);
  wire tmp6510;
  assign tmp6510 = 1'b0;
  wire tmp6511;
  assign tmp6511 = 1'b0;
  wire tmp6512;
  assign tmp6512 = 1'b0;
  wire tmp6513;
  assign tmp6513 = (tmp6510 & tmp6511) | (tmp6510 & tmp6512) | (tmp6511 & tmp6512);
  wire tmp6514;
  assign tmp6514 = (tmp6505 & tmp6509) | (tmp6505 & tmp6513) | (tmp6509 & tmp6513);
  wire tmp6515;
  assign tmp6515 = (tmp6488 & tmp6501) | (tmp6488 & tmp6514) | (tmp6501 & tmp6514);
  wire tmp6516;
  assign tmp6516 = 1'b0;
  wire tmp6517;
  assign tmp6517 = 1'b0;
  wire tmp6518;
  assign tmp6518 = 1'b0;
  wire tmp6519;
  assign tmp6519 = (tmp6516 & tmp6517) | (tmp6516 & tmp6518) | (tmp6517 & tmp6518);
  wire tmp6520;
  assign tmp6520 = 1'b0;
  wire tmp6521;
  assign tmp6521 = 1'b0;
  wire tmp6522;
  assign tmp6522 = 1'b0;
  wire tmp6523;
  assign tmp6523 = (tmp6520 & tmp6521) | (tmp6520 & tmp6522) | (tmp6521 & tmp6522);
  wire tmp6524;
  assign tmp6524 = 1'b0;
  wire tmp6525;
  assign tmp6525 = 1'b0;
  wire tmp6526;
  assign tmp6526 = 1'b0;
  wire tmp6527;
  assign tmp6527 = (tmp6524 & tmp6525) | (tmp6524 & tmp6526) | (tmp6525 & tmp6526);
  wire tmp6528;
  assign tmp6528 = (tmp6519 & tmp6523) | (tmp6519 & tmp6527) | (tmp6523 & tmp6527);
  wire tmp6529;
  assign tmp6529 = 1'b0;
  wire tmp6530;
  assign tmp6530 = 1'b0;
  wire tmp6531;
  assign tmp6531 = 1'b0;
  wire tmp6532;
  assign tmp6532 = (tmp6529 & tmp6530) | (tmp6529 & tmp6531) | (tmp6530 & tmp6531);
  wire tmp6533;
  assign tmp6533 = 1'b0;
  wire tmp6534;
  assign tmp6534 = 1'b0;
  wire tmp6535;
  assign tmp6535 = 1'b0;
  wire tmp6536;
  assign tmp6536 = (tmp6533 & tmp6534) | (tmp6533 & tmp6535) | (tmp6534 & tmp6535);
  wire tmp6537;
  assign tmp6537 = 1'b0;
  wire tmp6538;
  assign tmp6538 = 1'b0;
  wire tmp6539;
  assign tmp6539 = 1'b0;
  wire tmp6540;
  assign tmp6540 = (tmp6537 & tmp6538) | (tmp6537 & tmp6539) | (tmp6538 & tmp6539);
  wire tmp6541;
  assign tmp6541 = (tmp6532 & tmp6536) | (tmp6532 & tmp6540) | (tmp6536 & tmp6540);
  wire tmp6542;
  assign tmp6542 = 1'b0;
  wire tmp6543;
  assign tmp6543 = 1'b0;
  wire tmp6544;
  assign tmp6544 = 1'b0;
  wire tmp6545;
  assign tmp6545 = (tmp6542 & tmp6543) | (tmp6542 & tmp6544) | (tmp6543 & tmp6544);
  wire tmp6546;
  assign tmp6546 = 1'b0;
  wire tmp6547;
  assign tmp6547 = 1'b0;
  wire tmp6548;
  assign tmp6548 = 1'b0;
  wire tmp6549;
  assign tmp6549 = (tmp6546 & tmp6547) | (tmp6546 & tmp6548) | (tmp6547 & tmp6548);
  wire tmp6550;
  assign tmp6550 = 1'b0;
  wire tmp6551;
  assign tmp6551 = 1'b0;
  wire tmp6552;
  assign tmp6552 = 1'b0;
  wire tmp6553;
  assign tmp6553 = (tmp6550 & tmp6551) | (tmp6550 & tmp6552) | (tmp6551 & tmp6552);
  wire tmp6554;
  assign tmp6554 = (tmp6545 & tmp6549) | (tmp6545 & tmp6553) | (tmp6549 & tmp6553);
  wire tmp6555;
  assign tmp6555 = (tmp6528 & tmp6541) | (tmp6528 & tmp6554) | (tmp6541 & tmp6554);
  wire tmp6556;
  assign tmp6556 = (tmp6475 & tmp6515) | (tmp6475 & tmp6555) | (tmp6515 & tmp6555);
  wire tmp6557;
  assign tmp6557 = (tmp6314 & tmp6435) | (tmp6314 & tmp6556) | (tmp6435 & tmp6556);
  wire tmp6558;
  assign tmp6558 = (tmp5829 & tmp6193) | (tmp5829 & tmp6557) | (tmp6193 & tmp6557);
  wire tmp6559;
  assign tmp6559 = (tmp4372 & tmp5465) | (tmp4372 & tmp6558) | (tmp5465 & tmp6558);
  wire tmp6560;
  assign tmp6560 = 1'b0;
  wire tmp6561;
  assign tmp6561 = 1'b0;
  wire tmp6562;
  assign tmp6562 = 1'b0;
  wire tmp6563;
  assign tmp6563 = (tmp6560 & tmp6561) | (tmp6560 & tmp6562) | (tmp6561 & tmp6562);
  wire tmp6564;
  assign tmp6564 = 1'b0;
  wire tmp6565;
  assign tmp6565 = 1'b0;
  wire tmp6566;
  assign tmp6566 = 1'b0;
  wire tmp6567;
  assign tmp6567 = (tmp6564 & tmp6565) | (tmp6564 & tmp6566) | (tmp6565 & tmp6566);
  wire tmp6568;
  assign tmp6568 = 1'b0;
  wire tmp6569;
  assign tmp6569 = 1'b0;
  wire tmp6570;
  assign tmp6570 = 1'b0;
  wire tmp6571;
  assign tmp6571 = (tmp6568 & tmp6569) | (tmp6568 & tmp6570) | (tmp6569 & tmp6570);
  wire tmp6572;
  assign tmp6572 = (tmp6563 & tmp6567) | (tmp6563 & tmp6571) | (tmp6567 & tmp6571);
  wire tmp6573;
  assign tmp6573 = 1'b0;
  wire tmp6574;
  assign tmp6574 = 1'b0;
  wire tmp6575;
  assign tmp6575 = 1'b0;
  wire tmp6576;
  assign tmp6576 = (tmp6573 & tmp6574) | (tmp6573 & tmp6575) | (tmp6574 & tmp6575);
  wire tmp6577;
  assign tmp6577 = 1'b0;
  wire tmp6578;
  assign tmp6578 = 1'b0;
  wire tmp6579;
  assign tmp6579 = 1'b0;
  wire tmp6580;
  assign tmp6580 = (tmp6577 & tmp6578) | (tmp6577 & tmp6579) | (tmp6578 & tmp6579);
  wire tmp6581;
  assign tmp6581 = 1'b0;
  wire tmp6582;
  assign tmp6582 = 1'b0;
  wire tmp6583;
  assign tmp6583 = 1'b0;
  wire tmp6584;
  assign tmp6584 = (tmp6581 & tmp6582) | (tmp6581 & tmp6583) | (tmp6582 & tmp6583);
  wire tmp6585;
  assign tmp6585 = (tmp6576 & tmp6580) | (tmp6576 & tmp6584) | (tmp6580 & tmp6584);
  wire tmp6586;
  assign tmp6586 = 1'b0;
  wire tmp6587;
  assign tmp6587 = 1'b0;
  wire tmp6588;
  assign tmp6588 = 1'b0;
  wire tmp6589;
  assign tmp6589 = (tmp6586 & tmp6587) | (tmp6586 & tmp6588) | (tmp6587 & tmp6588);
  wire tmp6590;
  assign tmp6590 = 1'b0;
  wire tmp6591;
  assign tmp6591 = 1'b0;
  wire tmp6592;
  assign tmp6592 = 1'b0;
  wire tmp6593;
  assign tmp6593 = (tmp6590 & tmp6591) | (tmp6590 & tmp6592) | (tmp6591 & tmp6592);
  wire tmp6594;
  assign tmp6594 = 1'b0;
  wire tmp6595;
  assign tmp6595 = 1'b0;
  wire tmp6596;
  assign tmp6596 = 1'b0;
  wire tmp6597;
  assign tmp6597 = (tmp6594 & tmp6595) | (tmp6594 & tmp6596) | (tmp6595 & tmp6596);
  wire tmp6598;
  assign tmp6598 = (tmp6589 & tmp6593) | (tmp6589 & tmp6597) | (tmp6593 & tmp6597);
  wire tmp6599;
  assign tmp6599 = (tmp6572 & tmp6585) | (tmp6572 & tmp6598) | (tmp6585 & tmp6598);
  wire tmp6600;
  assign tmp6600 = 1'b0;
  wire tmp6601;
  assign tmp6601 = 1'b0;
  wire tmp6602;
  assign tmp6602 = 1'b0;
  wire tmp6603;
  assign tmp6603 = (tmp6600 & tmp6601) | (tmp6600 & tmp6602) | (tmp6601 & tmp6602);
  wire tmp6604;
  assign tmp6604 = 1'b0;
  wire tmp6605;
  assign tmp6605 = 1'b0;
  wire tmp6606;
  assign tmp6606 = 1'b0;
  wire tmp6607;
  assign tmp6607 = (tmp6604 & tmp6605) | (tmp6604 & tmp6606) | (tmp6605 & tmp6606);
  wire tmp6608;
  assign tmp6608 = 1'b0;
  wire tmp6609;
  assign tmp6609 = 1'b0;
  wire tmp6610;
  assign tmp6610 = 1'b0;
  wire tmp6611;
  assign tmp6611 = (tmp6608 & tmp6609) | (tmp6608 & tmp6610) | (tmp6609 & tmp6610);
  wire tmp6612;
  assign tmp6612 = (tmp6603 & tmp6607) | (tmp6603 & tmp6611) | (tmp6607 & tmp6611);
  wire tmp6613;
  assign tmp6613 = 1'b0;
  wire tmp6614;
  assign tmp6614 = 1'b0;
  wire tmp6615;
  assign tmp6615 = 1'b0;
  wire tmp6616;
  assign tmp6616 = (tmp6613 & tmp6614) | (tmp6613 & tmp6615) | (tmp6614 & tmp6615);
  wire tmp6617;
  assign tmp6617 = 1'b0;
  wire tmp6618;
  assign tmp6618 = 1'b1;
  wire tmp6619;
  assign tmp6619 = 1'b0;
  wire tmp6620;
  assign tmp6620 = (tmp6617 & tmp6618) | (tmp6617 & tmp6619) | (tmp6618 & tmp6619);
  wire tmp6621;
  assign tmp6621 = 1'b0;
  wire tmp6622;
  assign tmp6622 = 1'b0;
  wire tmp6623;
  assign tmp6623 = 1'b0;
  wire tmp6624;
  assign tmp6624 = (tmp6621 & tmp6622) | (tmp6621 & tmp6623) | (tmp6622 & tmp6623);
  wire tmp6625;
  assign tmp6625 = (tmp6616 & tmp6620) | (tmp6616 & tmp6624) | (tmp6620 & tmp6624);
  wire tmp6626;
  assign tmp6626 = 1'b0;
  wire tmp6627;
  assign tmp6627 = 1'b0;
  wire tmp6628;
  assign tmp6628 = 1'b0;
  wire tmp6629;
  assign tmp6629 = (tmp6626 & tmp6627) | (tmp6626 & tmp6628) | (tmp6627 & tmp6628);
  wire tmp6630;
  assign tmp6630 = 1'b0;
  wire tmp6631;
  assign tmp6631 = 1'b0;
  wire tmp6632;
  assign tmp6632 = 1'b0;
  wire tmp6633;
  assign tmp6633 = (tmp6630 & tmp6631) | (tmp6630 & tmp6632) | (tmp6631 & tmp6632);
  wire tmp6634;
  assign tmp6634 = 1'b0;
  wire tmp6635;
  assign tmp6635 = 1'b0;
  wire tmp6636;
  assign tmp6636 = 1'b0;
  wire tmp6637;
  assign tmp6637 = (tmp6634 & tmp6635) | (tmp6634 & tmp6636) | (tmp6635 & tmp6636);
  wire tmp6638;
  assign tmp6638 = (tmp6629 & tmp6633) | (tmp6629 & tmp6637) | (tmp6633 & tmp6637);
  wire tmp6639;
  assign tmp6639 = (tmp6612 & tmp6625) | (tmp6612 & tmp6638) | (tmp6625 & tmp6638);
  wire tmp6640;
  assign tmp6640 = 1'b0;
  wire tmp6641;
  assign tmp6641 = 1'b0;
  wire tmp6642;
  assign tmp6642 = 1'b0;
  wire tmp6643;
  assign tmp6643 = (tmp6640 & tmp6641) | (tmp6640 & tmp6642) | (tmp6641 & tmp6642);
  wire tmp6644;
  assign tmp6644 = 1'b0;
  wire tmp6645;
  assign tmp6645 = 1'b0;
  wire tmp6646;
  assign tmp6646 = 1'b0;
  wire tmp6647;
  assign tmp6647 = (tmp6644 & tmp6645) | (tmp6644 & tmp6646) | (tmp6645 & tmp6646);
  wire tmp6648;
  assign tmp6648 = 1'b0;
  wire tmp6649;
  assign tmp6649 = 1'b0;
  wire tmp6650;
  assign tmp6650 = 1'b0;
  wire tmp6651;
  assign tmp6651 = (tmp6648 & tmp6649) | (tmp6648 & tmp6650) | (tmp6649 & tmp6650);
  wire tmp6652;
  assign tmp6652 = (tmp6643 & tmp6647) | (tmp6643 & tmp6651) | (tmp6647 & tmp6651);
  wire tmp6653;
  assign tmp6653 = 1'b0;
  wire tmp6654;
  assign tmp6654 = 1'b0;
  wire tmp6655;
  assign tmp6655 = 1'b0;
  wire tmp6656;
  assign tmp6656 = (tmp6653 & tmp6654) | (tmp6653 & tmp6655) | (tmp6654 & tmp6655);
  wire tmp6657;
  assign tmp6657 = 1'b0;
  wire tmp6658;
  assign tmp6658 = 1'b0;
  wire tmp6659;
  assign tmp6659 = 1'b0;
  wire tmp6660;
  assign tmp6660 = (tmp6657 & tmp6658) | (tmp6657 & tmp6659) | (tmp6658 & tmp6659);
  wire tmp6661;
  assign tmp6661 = 1'b0;
  wire tmp6662;
  assign tmp6662 = 1'b0;
  wire tmp6663;
  assign tmp6663 = 1'b0;
  wire tmp6664;
  assign tmp6664 = (tmp6661 & tmp6662) | (tmp6661 & tmp6663) | (tmp6662 & tmp6663);
  wire tmp6665;
  assign tmp6665 = (tmp6656 & tmp6660) | (tmp6656 & tmp6664) | (tmp6660 & tmp6664);
  wire tmp6666;
  assign tmp6666 = 1'b0;
  wire tmp6667;
  assign tmp6667 = 1'b0;
  wire tmp6668;
  assign tmp6668 = 1'b0;
  wire tmp6669;
  assign tmp6669 = (tmp6666 & tmp6667) | (tmp6666 & tmp6668) | (tmp6667 & tmp6668);
  wire tmp6670;
  assign tmp6670 = 1'b0;
  wire tmp6671;
  assign tmp6671 = 1'b0;
  wire tmp6672;
  assign tmp6672 = 1'b0;
  wire tmp6673;
  assign tmp6673 = (tmp6670 & tmp6671) | (tmp6670 & tmp6672) | (tmp6671 & tmp6672);
  wire tmp6674;
  assign tmp6674 = 1'b0;
  wire tmp6675;
  assign tmp6675 = 1'b0;
  wire tmp6676;
  assign tmp6676 = 1'b0;
  wire tmp6677;
  assign tmp6677 = (tmp6674 & tmp6675) | (tmp6674 & tmp6676) | (tmp6675 & tmp6676);
  wire tmp6678;
  assign tmp6678 = (tmp6669 & tmp6673) | (tmp6669 & tmp6677) | (tmp6673 & tmp6677);
  wire tmp6679;
  assign tmp6679 = (tmp6652 & tmp6665) | (tmp6652 & tmp6678) | (tmp6665 & tmp6678);
  wire tmp6680;
  assign tmp6680 = (tmp6599 & tmp6639) | (tmp6599 & tmp6679) | (tmp6639 & tmp6679);
  wire tmp6681;
  assign tmp6681 = 1'b0;
  wire tmp6682;
  assign tmp6682 = 1'b0;
  wire tmp6683;
  assign tmp6683 = 1'b0;
  wire tmp6684;
  assign tmp6684 = (tmp6681 & tmp6682) | (tmp6681 & tmp6683) | (tmp6682 & tmp6683);
  wire tmp6685;
  assign tmp6685 = 1'b0;
  wire tmp6686;
  assign tmp6686 = 1'b0;
  wire tmp6687;
  assign tmp6687 = 1'b0;
  wire tmp6688;
  assign tmp6688 = (tmp6685 & tmp6686) | (tmp6685 & tmp6687) | (tmp6686 & tmp6687);
  wire tmp6689;
  assign tmp6689 = 1'b0;
  wire tmp6690;
  assign tmp6690 = 1'b0;
  wire tmp6691;
  assign tmp6691 = 1'b0;
  wire tmp6692;
  assign tmp6692 = (tmp6689 & tmp6690) | (tmp6689 & tmp6691) | (tmp6690 & tmp6691);
  wire tmp6693;
  assign tmp6693 = (tmp6684 & tmp6688) | (tmp6684 & tmp6692) | (tmp6688 & tmp6692);
  wire tmp6694;
  assign tmp6694 = 1'b0;
  wire tmp6695;
  assign tmp6695 = 1'b0;
  wire tmp6696;
  assign tmp6696 = 1'b0;
  wire tmp6697;
  assign tmp6697 = (tmp6694 & tmp6695) | (tmp6694 & tmp6696) | (tmp6695 & tmp6696);
  wire tmp6698;
  assign tmp6698 = 1'b0;
  wire tmp6699;
  assign tmp6699 = 1'b1;
  wire tmp6700;
  assign tmp6700 = 1'b0;
  wire tmp6701;
  assign tmp6701 = (tmp6698 & tmp6699) | (tmp6698 & tmp6700) | (tmp6699 & tmp6700);
  wire tmp6702;
  assign tmp6702 = 1'b0;
  wire tmp6703;
  assign tmp6703 = 1'b0;
  wire tmp6704;
  assign tmp6704 = 1'b0;
  wire tmp6705;
  assign tmp6705 = (tmp6702 & tmp6703) | (tmp6702 & tmp6704) | (tmp6703 & tmp6704);
  wire tmp6706;
  assign tmp6706 = (tmp6697 & tmp6701) | (tmp6697 & tmp6705) | (tmp6701 & tmp6705);
  wire tmp6707;
  assign tmp6707 = 1'b0;
  wire tmp6708;
  assign tmp6708 = 1'b0;
  wire tmp6709;
  assign tmp6709 = 1'b0;
  wire tmp6710;
  assign tmp6710 = (tmp6707 & tmp6708) | (tmp6707 & tmp6709) | (tmp6708 & tmp6709);
  wire tmp6711;
  assign tmp6711 = 1'b0;
  wire tmp6712;
  assign tmp6712 = 1'b0;
  wire tmp6713;
  assign tmp6713 = 1'b0;
  wire tmp6714;
  assign tmp6714 = (tmp6711 & tmp6712) | (tmp6711 & tmp6713) | (tmp6712 & tmp6713);
  wire tmp6715;
  assign tmp6715 = 1'b0;
  wire tmp6716;
  assign tmp6716 = 1'b0;
  wire tmp6717;
  assign tmp6717 = 1'b0;
  wire tmp6718;
  assign tmp6718 = (tmp6715 & tmp6716) | (tmp6715 & tmp6717) | (tmp6716 & tmp6717);
  wire tmp6719;
  assign tmp6719 = (tmp6710 & tmp6714) | (tmp6710 & tmp6718) | (tmp6714 & tmp6718);
  wire tmp6720;
  assign tmp6720 = (tmp6693 & tmp6706) | (tmp6693 & tmp6719) | (tmp6706 & tmp6719);
  wire tmp6721;
  assign tmp6721 = 1'b0;
  wire tmp6722;
  assign tmp6722 = 1'b0;
  wire tmp6723;
  assign tmp6723 = 1'b0;
  wire tmp6724;
  assign tmp6724 = (tmp6721 & tmp6722) | (tmp6721 & tmp6723) | (tmp6722 & tmp6723);
  wire tmp6725;
  assign tmp6725 = 1'b0;
  wire tmp6726;
  assign tmp6726 = 1'b1;
  wire tmp6727;
  assign tmp6727 = 1'b0;
  wire tmp6728;
  assign tmp6728 = (tmp6725 & tmp6726) | (tmp6725 & tmp6727) | (tmp6726 & tmp6727);
  wire tmp6729;
  assign tmp6729 = 1'b0;
  wire tmp6730;
  assign tmp6730 = 1'b0;
  wire tmp6731;
  assign tmp6731 = 1'b0;
  wire tmp6732;
  assign tmp6732 = (tmp6729 & tmp6730) | (tmp6729 & tmp6731) | (tmp6730 & tmp6731);
  wire tmp6733;
  assign tmp6733 = (tmp6724 & tmp6728) | (tmp6724 & tmp6732) | (tmp6728 & tmp6732);
  wire tmp6734;
  assign tmp6734 = 1'b0;
  wire tmp6735;
  assign tmp6735 = 1'b1;
  wire tmp6736;
  assign tmp6736 = 1'b0;
  wire tmp6737;
  assign tmp6737 = (tmp6734 & tmp6735) | (tmp6734 & tmp6736) | (tmp6735 & tmp6736);
  wire tmp6738;
  assign tmp6738 = 1'b1;
  wire tmp6739;
  assign tmp6739 = 1'b1;
  wire tmp6740;
  assign tmp6740 = 1'b1;
  wire tmp6741;
  assign tmp6741 = (tmp6738 & tmp6739) | (tmp6738 & tmp6740) | (tmp6739 & tmp6740);
  wire tmp6742;
  assign tmp6742 = 1'b0;
  wire tmp6743;
  assign tmp6743 = 1'b1;
  wire tmp6744;
  assign tmp6744 = 1'b0;
  wire tmp6745;
  assign tmp6745 = (tmp6742 & tmp6743) | (tmp6742 & tmp6744) | (tmp6743 & tmp6744);
  wire tmp6746;
  assign tmp6746 = (tmp6737 & tmp6741) | (tmp6737 & tmp6745) | (tmp6741 & tmp6745);
  wire tmp6747;
  assign tmp6747 = 1'b0;
  wire tmp6748;
  assign tmp6748 = 1'b0;
  wire tmp6749;
  assign tmp6749 = 1'b0;
  wire tmp6750;
  assign tmp6750 = (tmp6747 & tmp6748) | (tmp6747 & tmp6749) | (tmp6748 & tmp6749);
  wire tmp6751;
  assign tmp6751 = 1'b0;
  wire tmp6752;
  assign tmp6752 = 1'b1;
  wire tmp6753;
  assign tmp6753 = 1'b0;
  wire tmp6754;
  assign tmp6754 = (tmp6751 & tmp6752) | (tmp6751 & tmp6753) | (tmp6752 & tmp6753);
  wire tmp6755;
  assign tmp6755 = 1'b0;
  wire tmp6756;
  assign tmp6756 = 1'b0;
  wire tmp6757;
  assign tmp6757 = 1'b0;
  wire tmp6758;
  assign tmp6758 = (tmp6755 & tmp6756) | (tmp6755 & tmp6757) | (tmp6756 & tmp6757);
  wire tmp6759;
  assign tmp6759 = (tmp6750 & tmp6754) | (tmp6750 & tmp6758) | (tmp6754 & tmp6758);
  wire tmp6760;
  assign tmp6760 = (tmp6733 & tmp6746) | (tmp6733 & tmp6759) | (tmp6746 & tmp6759);
  wire tmp6761;
  assign tmp6761 = 1'b0;
  wire tmp6762;
  assign tmp6762 = 1'b0;
  wire tmp6763;
  assign tmp6763 = 1'b0;
  wire tmp6764;
  assign tmp6764 = (tmp6761 & tmp6762) | (tmp6761 & tmp6763) | (tmp6762 & tmp6763);
  wire tmp6765;
  assign tmp6765 = 1'b0;
  wire tmp6766;
  assign tmp6766 = 1'b0;
  wire tmp6767;
  assign tmp6767 = 1'b0;
  wire tmp6768;
  assign tmp6768 = (tmp6765 & tmp6766) | (tmp6765 & tmp6767) | (tmp6766 & tmp6767);
  wire tmp6769;
  assign tmp6769 = 1'b0;
  wire tmp6770;
  assign tmp6770 = 1'b0;
  wire tmp6771;
  assign tmp6771 = 1'b0;
  wire tmp6772;
  assign tmp6772 = (tmp6769 & tmp6770) | (tmp6769 & tmp6771) | (tmp6770 & tmp6771);
  wire tmp6773;
  assign tmp6773 = (tmp6764 & tmp6768) | (tmp6764 & tmp6772) | (tmp6768 & tmp6772);
  wire tmp6774;
  assign tmp6774 = 1'b0;
  wire tmp6775;
  assign tmp6775 = 1'b0;
  wire tmp6776;
  assign tmp6776 = 1'b0;
  wire tmp6777;
  assign tmp6777 = (tmp6774 & tmp6775) | (tmp6774 & tmp6776) | (tmp6775 & tmp6776);
  wire tmp6778;
  assign tmp6778 = 1'b0;
  wire tmp6779;
  assign tmp6779 = 1'b1;
  wire tmp6780;
  assign tmp6780 = 1'b0;
  wire tmp6781;
  assign tmp6781 = (tmp6778 & tmp6779) | (tmp6778 & tmp6780) | (tmp6779 & tmp6780);
  wire tmp6782;
  assign tmp6782 = 1'b0;
  wire tmp6783;
  assign tmp6783 = 1'b0;
  wire tmp6784;
  assign tmp6784 = 1'b0;
  wire tmp6785;
  assign tmp6785 = (tmp6782 & tmp6783) | (tmp6782 & tmp6784) | (tmp6783 & tmp6784);
  wire tmp6786;
  assign tmp6786 = (tmp6777 & tmp6781) | (tmp6777 & tmp6785) | (tmp6781 & tmp6785);
  wire tmp6787;
  assign tmp6787 = 1'b0;
  wire tmp6788;
  assign tmp6788 = 1'b0;
  wire tmp6789;
  assign tmp6789 = 1'b0;
  wire tmp6790;
  assign tmp6790 = (tmp6787 & tmp6788) | (tmp6787 & tmp6789) | (tmp6788 & tmp6789);
  wire tmp6791;
  assign tmp6791 = 1'b0;
  wire tmp6792;
  assign tmp6792 = 1'b0;
  wire tmp6793;
  assign tmp6793 = 1'b0;
  wire tmp6794;
  assign tmp6794 = (tmp6791 & tmp6792) | (tmp6791 & tmp6793) | (tmp6792 & tmp6793);
  wire tmp6795;
  assign tmp6795 = 1'b0;
  wire tmp6796;
  assign tmp6796 = 1'b0;
  wire tmp6797;
  assign tmp6797 = 1'b0;
  wire tmp6798;
  assign tmp6798 = (tmp6795 & tmp6796) | (tmp6795 & tmp6797) | (tmp6796 & tmp6797);
  wire tmp6799;
  assign tmp6799 = (tmp6790 & tmp6794) | (tmp6790 & tmp6798) | (tmp6794 & tmp6798);
  wire tmp6800;
  assign tmp6800 = (tmp6773 & tmp6786) | (tmp6773 & tmp6799) | (tmp6786 & tmp6799);
  wire tmp6801;
  assign tmp6801 = (tmp6720 & tmp6760) | (tmp6720 & tmp6800) | (tmp6760 & tmp6800);
  wire tmp6802;
  assign tmp6802 = 1'b0;
  wire tmp6803;
  assign tmp6803 = 1'b0;
  wire tmp6804;
  assign tmp6804 = 1'b0;
  wire tmp6805;
  assign tmp6805 = (tmp6802 & tmp6803) | (tmp6802 & tmp6804) | (tmp6803 & tmp6804);
  wire tmp6806;
  assign tmp6806 = 1'b0;
  wire tmp6807;
  assign tmp6807 = 1'b0;
  wire tmp6808;
  assign tmp6808 = 1'b0;
  wire tmp6809;
  assign tmp6809 = (tmp6806 & tmp6807) | (tmp6806 & tmp6808) | (tmp6807 & tmp6808);
  wire tmp6810;
  assign tmp6810 = 1'b0;
  wire tmp6811;
  assign tmp6811 = 1'b0;
  wire tmp6812;
  assign tmp6812 = 1'b0;
  wire tmp6813;
  assign tmp6813 = (tmp6810 & tmp6811) | (tmp6810 & tmp6812) | (tmp6811 & tmp6812);
  wire tmp6814;
  assign tmp6814 = (tmp6805 & tmp6809) | (tmp6805 & tmp6813) | (tmp6809 & tmp6813);
  wire tmp6815;
  assign tmp6815 = 1'b0;
  wire tmp6816;
  assign tmp6816 = 1'b0;
  wire tmp6817;
  assign tmp6817 = 1'b0;
  wire tmp6818;
  assign tmp6818 = (tmp6815 & tmp6816) | (tmp6815 & tmp6817) | (tmp6816 & tmp6817);
  wire tmp6819;
  assign tmp6819 = 1'b0;
  wire tmp6820;
  assign tmp6820 = 1'b0;
  wire tmp6821;
  assign tmp6821 = 1'b0;
  wire tmp6822;
  assign tmp6822 = (tmp6819 & tmp6820) | (tmp6819 & tmp6821) | (tmp6820 & tmp6821);
  wire tmp6823;
  assign tmp6823 = 1'b0;
  wire tmp6824;
  assign tmp6824 = 1'b0;
  wire tmp6825;
  assign tmp6825 = 1'b0;
  wire tmp6826;
  assign tmp6826 = (tmp6823 & tmp6824) | (tmp6823 & tmp6825) | (tmp6824 & tmp6825);
  wire tmp6827;
  assign tmp6827 = (tmp6818 & tmp6822) | (tmp6818 & tmp6826) | (tmp6822 & tmp6826);
  wire tmp6828;
  assign tmp6828 = 1'b0;
  wire tmp6829;
  assign tmp6829 = 1'b0;
  wire tmp6830;
  assign tmp6830 = 1'b0;
  wire tmp6831;
  assign tmp6831 = (tmp6828 & tmp6829) | (tmp6828 & tmp6830) | (tmp6829 & tmp6830);
  wire tmp6832;
  assign tmp6832 = 1'b0;
  wire tmp6833;
  assign tmp6833 = 1'b0;
  wire tmp6834;
  assign tmp6834 = 1'b0;
  wire tmp6835;
  assign tmp6835 = (tmp6832 & tmp6833) | (tmp6832 & tmp6834) | (tmp6833 & tmp6834);
  wire tmp6836;
  assign tmp6836 = 1'b0;
  wire tmp6837;
  assign tmp6837 = 1'b0;
  wire tmp6838;
  assign tmp6838 = 1'b0;
  wire tmp6839;
  assign tmp6839 = (tmp6836 & tmp6837) | (tmp6836 & tmp6838) | (tmp6837 & tmp6838);
  wire tmp6840;
  assign tmp6840 = (tmp6831 & tmp6835) | (tmp6831 & tmp6839) | (tmp6835 & tmp6839);
  wire tmp6841;
  assign tmp6841 = (tmp6814 & tmp6827) | (tmp6814 & tmp6840) | (tmp6827 & tmp6840);
  wire tmp6842;
  assign tmp6842 = 1'b0;
  wire tmp6843;
  assign tmp6843 = 1'b0;
  wire tmp6844;
  assign tmp6844 = 1'b0;
  wire tmp6845;
  assign tmp6845 = (tmp6842 & tmp6843) | (tmp6842 & tmp6844) | (tmp6843 & tmp6844);
  wire tmp6846;
  assign tmp6846 = 1'b0;
  wire tmp6847;
  assign tmp6847 = 1'b0;
  wire tmp6848;
  assign tmp6848 = 1'b0;
  wire tmp6849;
  assign tmp6849 = (tmp6846 & tmp6847) | (tmp6846 & tmp6848) | (tmp6847 & tmp6848);
  wire tmp6850;
  assign tmp6850 = 1'b0;
  wire tmp6851;
  assign tmp6851 = 1'b0;
  wire tmp6852;
  assign tmp6852 = 1'b0;
  wire tmp6853;
  assign tmp6853 = (tmp6850 & tmp6851) | (tmp6850 & tmp6852) | (tmp6851 & tmp6852);
  wire tmp6854;
  assign tmp6854 = (tmp6845 & tmp6849) | (tmp6845 & tmp6853) | (tmp6849 & tmp6853);
  wire tmp6855;
  assign tmp6855 = 1'b0;
  wire tmp6856;
  assign tmp6856 = 1'b0;
  wire tmp6857;
  assign tmp6857 = 1'b0;
  wire tmp6858;
  assign tmp6858 = (tmp6855 & tmp6856) | (tmp6855 & tmp6857) | (tmp6856 & tmp6857);
  wire tmp6859;
  assign tmp6859 = 1'b0;
  wire tmp6860;
  assign tmp6860 = 1'b1;
  wire tmp6861;
  assign tmp6861 = 1'b0;
  wire tmp6862;
  assign tmp6862 = (tmp6859 & tmp6860) | (tmp6859 & tmp6861) | (tmp6860 & tmp6861);
  wire tmp6863;
  assign tmp6863 = 1'b0;
  wire tmp6864;
  assign tmp6864 = 1'b0;
  wire tmp6865;
  assign tmp6865 = 1'b0;
  wire tmp6866;
  assign tmp6866 = (tmp6863 & tmp6864) | (tmp6863 & tmp6865) | (tmp6864 & tmp6865);
  wire tmp6867;
  assign tmp6867 = (tmp6858 & tmp6862) | (tmp6858 & tmp6866) | (tmp6862 & tmp6866);
  wire tmp6868;
  assign tmp6868 = 1'b0;
  wire tmp6869;
  assign tmp6869 = 1'b0;
  wire tmp6870;
  assign tmp6870 = 1'b0;
  wire tmp6871;
  assign tmp6871 = (tmp6868 & tmp6869) | (tmp6868 & tmp6870) | (tmp6869 & tmp6870);
  wire tmp6872;
  assign tmp6872 = 1'b0;
  wire tmp6873;
  assign tmp6873 = 1'b0;
  wire tmp6874;
  assign tmp6874 = 1'b0;
  wire tmp6875;
  assign tmp6875 = (tmp6872 & tmp6873) | (tmp6872 & tmp6874) | (tmp6873 & tmp6874);
  wire tmp6876;
  assign tmp6876 = 1'b0;
  wire tmp6877;
  assign tmp6877 = 1'b0;
  wire tmp6878;
  assign tmp6878 = 1'b0;
  wire tmp6879;
  assign tmp6879 = (tmp6876 & tmp6877) | (tmp6876 & tmp6878) | (tmp6877 & tmp6878);
  wire tmp6880;
  assign tmp6880 = (tmp6871 & tmp6875) | (tmp6871 & tmp6879) | (tmp6875 & tmp6879);
  wire tmp6881;
  assign tmp6881 = (tmp6854 & tmp6867) | (tmp6854 & tmp6880) | (tmp6867 & tmp6880);
  wire tmp6882;
  assign tmp6882 = 1'b0;
  wire tmp6883;
  assign tmp6883 = 1'b0;
  wire tmp6884;
  assign tmp6884 = 1'b0;
  wire tmp6885;
  assign tmp6885 = (tmp6882 & tmp6883) | (tmp6882 & tmp6884) | (tmp6883 & tmp6884);
  wire tmp6886;
  assign tmp6886 = 1'b0;
  wire tmp6887;
  assign tmp6887 = 1'b0;
  wire tmp6888;
  assign tmp6888 = 1'b0;
  wire tmp6889;
  assign tmp6889 = (tmp6886 & tmp6887) | (tmp6886 & tmp6888) | (tmp6887 & tmp6888);
  wire tmp6890;
  assign tmp6890 = 1'b0;
  wire tmp6891;
  assign tmp6891 = 1'b0;
  wire tmp6892;
  assign tmp6892 = 1'b0;
  wire tmp6893;
  assign tmp6893 = (tmp6890 & tmp6891) | (tmp6890 & tmp6892) | (tmp6891 & tmp6892);
  wire tmp6894;
  assign tmp6894 = (tmp6885 & tmp6889) | (tmp6885 & tmp6893) | (tmp6889 & tmp6893);
  wire tmp6895;
  assign tmp6895 = 1'b0;
  wire tmp6896;
  assign tmp6896 = 1'b0;
  wire tmp6897;
  assign tmp6897 = 1'b0;
  wire tmp6898;
  assign tmp6898 = (tmp6895 & tmp6896) | (tmp6895 & tmp6897) | (tmp6896 & tmp6897);
  wire tmp6899;
  assign tmp6899 = 1'b0;
  wire tmp6900;
  assign tmp6900 = 1'b0;
  wire tmp6901;
  assign tmp6901 = 1'b0;
  wire tmp6902;
  assign tmp6902 = (tmp6899 & tmp6900) | (tmp6899 & tmp6901) | (tmp6900 & tmp6901);
  wire tmp6903;
  assign tmp6903 = 1'b0;
  wire tmp6904;
  assign tmp6904 = 1'b0;
  wire tmp6905;
  assign tmp6905 = 1'b0;
  wire tmp6906;
  assign tmp6906 = (tmp6903 & tmp6904) | (tmp6903 & tmp6905) | (tmp6904 & tmp6905);
  wire tmp6907;
  assign tmp6907 = (tmp6898 & tmp6902) | (tmp6898 & tmp6906) | (tmp6902 & tmp6906);
  wire tmp6908;
  assign tmp6908 = 1'b0;
  wire tmp6909;
  assign tmp6909 = 1'b0;
  wire tmp6910;
  assign tmp6910 = 1'b0;
  wire tmp6911;
  assign tmp6911 = (tmp6908 & tmp6909) | (tmp6908 & tmp6910) | (tmp6909 & tmp6910);
  wire tmp6912;
  assign tmp6912 = 1'b0;
  wire tmp6913;
  assign tmp6913 = 1'b0;
  wire tmp6914;
  assign tmp6914 = 1'b0;
  wire tmp6915;
  assign tmp6915 = (tmp6912 & tmp6913) | (tmp6912 & tmp6914) | (tmp6913 & tmp6914);
  wire tmp6916;
  assign tmp6916 = 1'b0;
  wire tmp6917;
  assign tmp6917 = 1'b0;
  wire tmp6918;
  assign tmp6918 = 1'b0;
  wire tmp6919;
  assign tmp6919 = (tmp6916 & tmp6917) | (tmp6916 & tmp6918) | (tmp6917 & tmp6918);
  wire tmp6920;
  assign tmp6920 = (tmp6911 & tmp6915) | (tmp6911 & tmp6919) | (tmp6915 & tmp6919);
  wire tmp6921;
  assign tmp6921 = (tmp6894 & tmp6907) | (tmp6894 & tmp6920) | (tmp6907 & tmp6920);
  wire tmp6922;
  assign tmp6922 = (tmp6841 & tmp6881) | (tmp6841 & tmp6921) | (tmp6881 & tmp6921);
  wire tmp6923;
  assign tmp6923 = (tmp6680 & tmp6801) | (tmp6680 & tmp6922) | (tmp6801 & tmp6922);
  wire tmp6924;
  assign tmp6924 = 1'b0;
  wire tmp6925;
  assign tmp6925 = 1'b0;
  wire tmp6926;
  assign tmp6926 = 1'b0;
  wire tmp6927;
  assign tmp6927 = (tmp6924 & tmp6925) | (tmp6924 & tmp6926) | (tmp6925 & tmp6926);
  wire tmp6928;
  assign tmp6928 = 1'b0;
  wire tmp6929;
  assign tmp6929 = 1'b0;
  wire tmp6930;
  assign tmp6930 = 1'b0;
  wire tmp6931;
  assign tmp6931 = (tmp6928 & tmp6929) | (tmp6928 & tmp6930) | (tmp6929 & tmp6930);
  wire tmp6932;
  assign tmp6932 = 1'b0;
  wire tmp6933;
  assign tmp6933 = 1'b0;
  wire tmp6934;
  assign tmp6934 = 1'b0;
  wire tmp6935;
  assign tmp6935 = (tmp6932 & tmp6933) | (tmp6932 & tmp6934) | (tmp6933 & tmp6934);
  wire tmp6936;
  assign tmp6936 = (tmp6927 & tmp6931) | (tmp6927 & tmp6935) | (tmp6931 & tmp6935);
  wire tmp6937;
  assign tmp6937 = 1'b0;
  wire tmp6938;
  assign tmp6938 = 1'b0;
  wire tmp6939;
  assign tmp6939 = 1'b0;
  wire tmp6940;
  assign tmp6940 = (tmp6937 & tmp6938) | (tmp6937 & tmp6939) | (tmp6938 & tmp6939);
  wire tmp6941;
  assign tmp6941 = 1'b0;
  wire tmp6942;
  assign tmp6942 = 1'b1;
  wire tmp6943;
  assign tmp6943 = 1'b0;
  wire tmp6944;
  assign tmp6944 = (tmp6941 & tmp6942) | (tmp6941 & tmp6943) | (tmp6942 & tmp6943);
  wire tmp6945;
  assign tmp6945 = 1'b0;
  wire tmp6946;
  assign tmp6946 = 1'b0;
  wire tmp6947;
  assign tmp6947 = 1'b0;
  wire tmp6948;
  assign tmp6948 = (tmp6945 & tmp6946) | (tmp6945 & tmp6947) | (tmp6946 & tmp6947);
  wire tmp6949;
  assign tmp6949 = (tmp6940 & tmp6944) | (tmp6940 & tmp6948) | (tmp6944 & tmp6948);
  wire tmp6950;
  assign tmp6950 = 1'b0;
  wire tmp6951;
  assign tmp6951 = 1'b0;
  wire tmp6952;
  assign tmp6952 = 1'b0;
  wire tmp6953;
  assign tmp6953 = (tmp6950 & tmp6951) | (tmp6950 & tmp6952) | (tmp6951 & tmp6952);
  wire tmp6954;
  assign tmp6954 = 1'b0;
  wire tmp6955;
  assign tmp6955 = 1'b0;
  wire tmp6956;
  assign tmp6956 = 1'b0;
  wire tmp6957;
  assign tmp6957 = (tmp6954 & tmp6955) | (tmp6954 & tmp6956) | (tmp6955 & tmp6956);
  wire tmp6958;
  assign tmp6958 = 1'b0;
  wire tmp6959;
  assign tmp6959 = 1'b0;
  wire tmp6960;
  assign tmp6960 = 1'b0;
  wire tmp6961;
  assign tmp6961 = (tmp6958 & tmp6959) | (tmp6958 & tmp6960) | (tmp6959 & tmp6960);
  wire tmp6962;
  assign tmp6962 = (tmp6953 & tmp6957) | (tmp6953 & tmp6961) | (tmp6957 & tmp6961);
  wire tmp6963;
  assign tmp6963 = (tmp6936 & tmp6949) | (tmp6936 & tmp6962) | (tmp6949 & tmp6962);
  wire tmp6964;
  assign tmp6964 = 1'b0;
  wire tmp6965;
  assign tmp6965 = 1'b0;
  wire tmp6966;
  assign tmp6966 = 1'b0;
  wire tmp6967;
  assign tmp6967 = (tmp6964 & tmp6965) | (tmp6964 & tmp6966) | (tmp6965 & tmp6966);
  wire tmp6968;
  assign tmp6968 = 1'b0;
  wire tmp6969;
  assign tmp6969 = 1'b1;
  wire tmp6970;
  assign tmp6970 = 1'b0;
  wire tmp6971;
  assign tmp6971 = (tmp6968 & tmp6969) | (tmp6968 & tmp6970) | (tmp6969 & tmp6970);
  wire tmp6972;
  assign tmp6972 = 1'b0;
  wire tmp6973;
  assign tmp6973 = 1'b0;
  wire tmp6974;
  assign tmp6974 = 1'b0;
  wire tmp6975;
  assign tmp6975 = (tmp6972 & tmp6973) | (tmp6972 & tmp6974) | (tmp6973 & tmp6974);
  wire tmp6976;
  assign tmp6976 = (tmp6967 & tmp6971) | (tmp6967 & tmp6975) | (tmp6971 & tmp6975);
  wire tmp6977;
  assign tmp6977 = 1'b0;
  wire tmp6978;
  assign tmp6978 = 1'b1;
  wire tmp6979;
  assign tmp6979 = 1'b0;
  wire tmp6980;
  assign tmp6980 = (tmp6977 & tmp6978) | (tmp6977 & tmp6979) | (tmp6978 & tmp6979);
  wire tmp6981;
  assign tmp6981 = 1'b1;
  wire tmp6982;
  assign tmp6982 = 1'b1;
  wire tmp6983;
  assign tmp6983 = 1'b1;
  wire tmp6984;
  assign tmp6984 = (tmp6981 & tmp6982) | (tmp6981 & tmp6983) | (tmp6982 & tmp6983);
  wire tmp6985;
  assign tmp6985 = 1'b0;
  wire tmp6986;
  assign tmp6986 = 1'b1;
  wire tmp6987;
  assign tmp6987 = 1'b0;
  wire tmp6988;
  assign tmp6988 = (tmp6985 & tmp6986) | (tmp6985 & tmp6987) | (tmp6986 & tmp6987);
  wire tmp6989;
  assign tmp6989 = (tmp6980 & tmp6984) | (tmp6980 & tmp6988) | (tmp6984 & tmp6988);
  wire tmp6990;
  assign tmp6990 = 1'b0;
  wire tmp6991;
  assign tmp6991 = 1'b0;
  wire tmp6992;
  assign tmp6992 = 1'b0;
  wire tmp6993;
  assign tmp6993 = (tmp6990 & tmp6991) | (tmp6990 & tmp6992) | (tmp6991 & tmp6992);
  wire tmp6994;
  assign tmp6994 = 1'b0;
  wire tmp6995;
  assign tmp6995 = 1'b1;
  wire tmp6996;
  assign tmp6996 = 1'b0;
  wire tmp6997;
  assign tmp6997 = (tmp6994 & tmp6995) | (tmp6994 & tmp6996) | (tmp6995 & tmp6996);
  wire tmp6998;
  assign tmp6998 = 1'b0;
  wire tmp6999;
  assign tmp6999 = 1'b0;
  wire tmp7000;
  assign tmp7000 = 1'b0;
  wire tmp7001;
  assign tmp7001 = (tmp6998 & tmp6999) | (tmp6998 & tmp7000) | (tmp6999 & tmp7000);
  wire tmp7002;
  assign tmp7002 = (tmp6993 & tmp6997) | (tmp6993 & tmp7001) | (tmp6997 & tmp7001);
  wire tmp7003;
  assign tmp7003 = (tmp6976 & tmp6989) | (tmp6976 & tmp7002) | (tmp6989 & tmp7002);
  wire tmp7004;
  assign tmp7004 = 1'b0;
  wire tmp7005;
  assign tmp7005 = 1'b0;
  wire tmp7006;
  assign tmp7006 = 1'b0;
  wire tmp7007;
  assign tmp7007 = (tmp7004 & tmp7005) | (tmp7004 & tmp7006) | (tmp7005 & tmp7006);
  wire tmp7008;
  assign tmp7008 = 1'b0;
  wire tmp7009;
  assign tmp7009 = 1'b0;
  wire tmp7010;
  assign tmp7010 = 1'b0;
  wire tmp7011;
  assign tmp7011 = (tmp7008 & tmp7009) | (tmp7008 & tmp7010) | (tmp7009 & tmp7010);
  wire tmp7012;
  assign tmp7012 = 1'b0;
  wire tmp7013;
  assign tmp7013 = 1'b0;
  wire tmp7014;
  assign tmp7014 = 1'b0;
  wire tmp7015;
  assign tmp7015 = (tmp7012 & tmp7013) | (tmp7012 & tmp7014) | (tmp7013 & tmp7014);
  wire tmp7016;
  assign tmp7016 = (tmp7007 & tmp7011) | (tmp7007 & tmp7015) | (tmp7011 & tmp7015);
  wire tmp7017;
  assign tmp7017 = 1'b0;
  wire tmp7018;
  assign tmp7018 = 1'b0;
  wire tmp7019;
  assign tmp7019 = 1'b0;
  wire tmp7020;
  assign tmp7020 = (tmp7017 & tmp7018) | (tmp7017 & tmp7019) | (tmp7018 & tmp7019);
  wire tmp7021;
  assign tmp7021 = 1'b0;
  wire tmp7022;
  assign tmp7022 = 1'b1;
  wire tmp7023;
  assign tmp7023 = 1'b0;
  wire tmp7024;
  assign tmp7024 = (tmp7021 & tmp7022) | (tmp7021 & tmp7023) | (tmp7022 & tmp7023);
  wire tmp7025;
  assign tmp7025 = 1'b0;
  wire tmp7026;
  assign tmp7026 = 1'b0;
  wire tmp7027;
  assign tmp7027 = 1'b0;
  wire tmp7028;
  assign tmp7028 = (tmp7025 & tmp7026) | (tmp7025 & tmp7027) | (tmp7026 & tmp7027);
  wire tmp7029;
  assign tmp7029 = (tmp7020 & tmp7024) | (tmp7020 & tmp7028) | (tmp7024 & tmp7028);
  wire tmp7030;
  assign tmp7030 = 1'b0;
  wire tmp7031;
  assign tmp7031 = 1'b0;
  wire tmp7032;
  assign tmp7032 = 1'b0;
  wire tmp7033;
  assign tmp7033 = (tmp7030 & tmp7031) | (tmp7030 & tmp7032) | (tmp7031 & tmp7032);
  wire tmp7034;
  assign tmp7034 = 1'b0;
  wire tmp7035;
  assign tmp7035 = 1'b0;
  wire tmp7036;
  assign tmp7036 = 1'b0;
  wire tmp7037;
  assign tmp7037 = (tmp7034 & tmp7035) | (tmp7034 & tmp7036) | (tmp7035 & tmp7036);
  wire tmp7038;
  assign tmp7038 = 1'b0;
  wire tmp7039;
  assign tmp7039 = 1'b0;
  wire tmp7040;
  assign tmp7040 = 1'b0;
  wire tmp7041;
  assign tmp7041 = (tmp7038 & tmp7039) | (tmp7038 & tmp7040) | (tmp7039 & tmp7040);
  wire tmp7042;
  assign tmp7042 = (tmp7033 & tmp7037) | (tmp7033 & tmp7041) | (tmp7037 & tmp7041);
  wire tmp7043;
  assign tmp7043 = (tmp7016 & tmp7029) | (tmp7016 & tmp7042) | (tmp7029 & tmp7042);
  wire tmp7044;
  assign tmp7044 = (tmp6963 & tmp7003) | (tmp6963 & tmp7043) | (tmp7003 & tmp7043);
  wire tmp7045;
  assign tmp7045 = 1'b0;
  wire tmp7046;
  assign tmp7046 = 1'b0;
  wire tmp7047;
  assign tmp7047 = 1'b0;
  wire tmp7048;
  assign tmp7048 = (tmp7045 & tmp7046) | (tmp7045 & tmp7047) | (tmp7046 & tmp7047);
  wire tmp7049;
  assign tmp7049 = 1'b0;
  wire tmp7050;
  assign tmp7050 = 1'b1;
  wire tmp7051;
  assign tmp7051 = 1'b0;
  wire tmp7052;
  assign tmp7052 = (tmp7049 & tmp7050) | (tmp7049 & tmp7051) | (tmp7050 & tmp7051);
  wire tmp7053;
  assign tmp7053 = 1'b0;
  wire tmp7054;
  assign tmp7054 = 1'b0;
  wire tmp7055;
  assign tmp7055 = 1'b0;
  wire tmp7056;
  assign tmp7056 = (tmp7053 & tmp7054) | (tmp7053 & tmp7055) | (tmp7054 & tmp7055);
  wire tmp7057;
  assign tmp7057 = (tmp7048 & tmp7052) | (tmp7048 & tmp7056) | (tmp7052 & tmp7056);
  wire tmp7058;
  assign tmp7058 = 1'b0;
  wire tmp7059;
  assign tmp7059 = 1'b1;
  wire tmp7060;
  assign tmp7060 = 1'b0;
  wire tmp7061;
  assign tmp7061 = (tmp7058 & tmp7059) | (tmp7058 & tmp7060) | (tmp7059 & tmp7060);
  wire tmp7062;
  assign tmp7062 = 1'b1;
  wire tmp7063;
  assign tmp7063 = 1'b1;
  wire tmp7064;
  assign tmp7064 = 1'b1;
  wire tmp7065;
  assign tmp7065 = (tmp7062 & tmp7063) | (tmp7062 & tmp7064) | (tmp7063 & tmp7064);
  wire tmp7066;
  assign tmp7066 = 1'b0;
  wire tmp7067;
  assign tmp7067 = 1'b1;
  wire tmp7068;
  assign tmp7068 = 1'b0;
  wire tmp7069;
  assign tmp7069 = (tmp7066 & tmp7067) | (tmp7066 & tmp7068) | (tmp7067 & tmp7068);
  wire tmp7070;
  assign tmp7070 = (tmp7061 & tmp7065) | (tmp7061 & tmp7069) | (tmp7065 & tmp7069);
  wire tmp7071;
  assign tmp7071 = 1'b0;
  wire tmp7072;
  assign tmp7072 = 1'b0;
  wire tmp7073;
  assign tmp7073 = 1'b0;
  wire tmp7074;
  assign tmp7074 = (tmp7071 & tmp7072) | (tmp7071 & tmp7073) | (tmp7072 & tmp7073);
  wire tmp7075;
  assign tmp7075 = 1'b0;
  wire tmp7076;
  assign tmp7076 = 1'b1;
  wire tmp7077;
  assign tmp7077 = 1'b0;
  wire tmp7078;
  assign tmp7078 = (tmp7075 & tmp7076) | (tmp7075 & tmp7077) | (tmp7076 & tmp7077);
  wire tmp7079;
  assign tmp7079 = 1'b0;
  wire tmp7080;
  assign tmp7080 = 1'b0;
  wire tmp7081;
  assign tmp7081 = 1'b0;
  wire tmp7082;
  assign tmp7082 = (tmp7079 & tmp7080) | (tmp7079 & tmp7081) | (tmp7080 & tmp7081);
  wire tmp7083;
  assign tmp7083 = (tmp7074 & tmp7078) | (tmp7074 & tmp7082) | (tmp7078 & tmp7082);
  wire tmp7084;
  assign tmp7084 = (tmp7057 & tmp7070) | (tmp7057 & tmp7083) | (tmp7070 & tmp7083);
  wire tmp7085;
  assign tmp7085 = 1'b0;
  wire tmp7086;
  assign tmp7086 = 1'b1;
  wire tmp7087;
  assign tmp7087 = 1'b0;
  wire tmp7088;
  assign tmp7088 = (tmp7085 & tmp7086) | (tmp7085 & tmp7087) | (tmp7086 & tmp7087);
  wire tmp7089;
  assign tmp7089 = 1'b1;
  wire tmp7090;
  assign tmp7090 = 1'b1;
  wire tmp7091;
  assign tmp7091 = 1'b1;
  wire tmp7092;
  assign tmp7092 = (tmp7089 & tmp7090) | (tmp7089 & tmp7091) | (tmp7090 & tmp7091);
  wire tmp7093;
  assign tmp7093 = 1'b0;
  wire tmp7094;
  assign tmp7094 = 1'b1;
  wire tmp7095;
  assign tmp7095 = 1'b0;
  wire tmp7096;
  assign tmp7096 = (tmp7093 & tmp7094) | (tmp7093 & tmp7095) | (tmp7094 & tmp7095);
  wire tmp7097;
  assign tmp7097 = (tmp7088 & tmp7092) | (tmp7088 & tmp7096) | (tmp7092 & tmp7096);
  wire tmp7098;
  assign tmp7098 = 1'b1;
  wire tmp7099;
  assign tmp7099 = 1'b1;
  wire tmp7100;
  assign tmp7100 = 1'b1;
  wire tmp7101;
  assign tmp7101 = (tmp7098 & tmp7099) | (tmp7098 & tmp7100) | (tmp7099 & tmp7100);
  wire tmp7102;
  assign tmp7102 = 1'b1;
  wire tmp7103;
  assign tmp7103 = ~pi5;
  wire tmp7104;
  assign tmp7104 = ~pi6;
  wire tmp7105;
  assign tmp7105 = (tmp7102 & tmp7103) | (tmp7102 & tmp7104) | (tmp7103 & tmp7104);
  wire tmp7106;
  assign tmp7106 = 1'b1;
  wire tmp7107;
  assign tmp7107 = ~pi6;
  wire tmp7108;
  assign tmp7108 = ~pi7;
  wire tmp7109;
  assign tmp7109 = (tmp7106 & tmp7107) | (tmp7106 & tmp7108) | (tmp7107 & tmp7108);
  wire tmp7110;
  assign tmp7110 = (tmp7101 & tmp7105) | (tmp7101 & tmp7109) | (tmp7105 & tmp7109);
  wire tmp7111;
  assign tmp7111 = 1'b0;
  wire tmp7112;
  assign tmp7112 = 1'b1;
  wire tmp7113;
  assign tmp7113 = 1'b0;
  wire tmp7114;
  assign tmp7114 = (tmp7111 & tmp7112) | (tmp7111 & tmp7113) | (tmp7112 & tmp7113);
  wire tmp7115;
  assign tmp7115 = 1'b1;
  wire tmp7116;
  assign tmp7116 = ~pi6;
  wire tmp7117;
  assign tmp7117 = ~pi7;
  wire tmp7118;
  assign tmp7118 = (tmp7115 & tmp7116) | (tmp7115 & tmp7117) | (tmp7116 & tmp7117);
  wire tmp7119;
  assign tmp7119 = 1'b0;
  wire tmp7120;
  assign tmp7120 = ~pi7;
  wire tmp7121;
  assign tmp7121 = 1'b0;
  wire tmp7122;
  assign tmp7122 = (tmp7119 & tmp7120) | (tmp7119 & tmp7121) | (tmp7120 & tmp7121);
  wire tmp7123;
  assign tmp7123 = (tmp7114 & tmp7118) | (tmp7114 & tmp7122) | (tmp7118 & tmp7122);
  wire tmp7124;
  assign tmp7124 = (tmp7097 & tmp7110) | (tmp7097 & tmp7123) | (tmp7110 & tmp7123);
  wire tmp7125;
  assign tmp7125 = 1'b0;
  wire tmp7126;
  assign tmp7126 = 1'b0;
  wire tmp7127;
  assign tmp7127 = 1'b0;
  wire tmp7128;
  assign tmp7128 = (tmp7125 & tmp7126) | (tmp7125 & tmp7127) | (tmp7126 & tmp7127);
  wire tmp7129;
  assign tmp7129 = 1'b0;
  wire tmp7130;
  assign tmp7130 = 1'b1;
  wire tmp7131;
  assign tmp7131 = 1'b0;
  wire tmp7132;
  assign tmp7132 = (tmp7129 & tmp7130) | (tmp7129 & tmp7131) | (tmp7130 & tmp7131);
  wire tmp7133;
  assign tmp7133 = 1'b0;
  wire tmp7134;
  assign tmp7134 = 1'b0;
  wire tmp7135;
  assign tmp7135 = 1'b0;
  wire tmp7136;
  assign tmp7136 = (tmp7133 & tmp7134) | (tmp7133 & tmp7135) | (tmp7134 & tmp7135);
  wire tmp7137;
  assign tmp7137 = (tmp7128 & tmp7132) | (tmp7128 & tmp7136) | (tmp7132 & tmp7136);
  wire tmp7138;
  assign tmp7138 = 1'b0;
  wire tmp7139;
  assign tmp7139 = 1'b1;
  wire tmp7140;
  assign tmp7140 = 1'b0;
  wire tmp7141;
  assign tmp7141 = (tmp7138 & tmp7139) | (tmp7138 & tmp7140) | (tmp7139 & tmp7140);
  wire tmp7142;
  assign tmp7142 = 1'b1;
  wire tmp7143;
  assign tmp7143 = ~pi6;
  wire tmp7144;
  assign tmp7144 = ~pi7;
  wire tmp7145;
  assign tmp7145 = (tmp7142 & tmp7143) | (tmp7142 & tmp7144) | (tmp7143 & tmp7144);
  wire tmp7146;
  assign tmp7146 = 1'b0;
  wire tmp7147;
  assign tmp7147 = ~pi7;
  wire tmp7148;
  assign tmp7148 = 1'b0;
  wire tmp7149;
  assign tmp7149 = (tmp7146 & tmp7147) | (tmp7146 & tmp7148) | (tmp7147 & tmp7148);
  wire tmp7150;
  assign tmp7150 = (tmp7141 & tmp7145) | (tmp7141 & tmp7149) | (tmp7145 & tmp7149);
  wire tmp7151;
  assign tmp7151 = 1'b0;
  wire tmp7152;
  assign tmp7152 = 1'b0;
  wire tmp7153;
  assign tmp7153 = 1'b0;
  wire tmp7154;
  assign tmp7154 = (tmp7151 & tmp7152) | (tmp7151 & tmp7153) | (tmp7152 & tmp7153);
  wire tmp7155;
  assign tmp7155 = 1'b0;
  wire tmp7156;
  assign tmp7156 = ~pi7;
  wire tmp7157;
  assign tmp7157 = 1'b0;
  wire tmp7158;
  assign tmp7158 = (tmp7155 & tmp7156) | (tmp7155 & tmp7157) | (tmp7156 & tmp7157);
  wire tmp7159;
  assign tmp7159 = 1'b0;
  wire tmp7160;
  assign tmp7160 = 1'b0;
  wire tmp7161;
  assign tmp7161 = 1'b0;
  wire tmp7162;
  assign tmp7162 = (tmp7159 & tmp7160) | (tmp7159 & tmp7161) | (tmp7160 & tmp7161);
  wire tmp7163;
  assign tmp7163 = (tmp7154 & tmp7158) | (tmp7154 & tmp7162) | (tmp7158 & tmp7162);
  wire tmp7164;
  assign tmp7164 = (tmp7137 & tmp7150) | (tmp7137 & tmp7163) | (tmp7150 & tmp7163);
  wire tmp7165;
  assign tmp7165 = (tmp7084 & tmp7124) | (tmp7084 & tmp7164) | (tmp7124 & tmp7164);
  wire tmp7166;
  assign tmp7166 = 1'b0;
  wire tmp7167;
  assign tmp7167 = 1'b0;
  wire tmp7168;
  assign tmp7168 = 1'b0;
  wire tmp7169;
  assign tmp7169 = (tmp7166 & tmp7167) | (tmp7166 & tmp7168) | (tmp7167 & tmp7168);
  wire tmp7170;
  assign tmp7170 = 1'b0;
  wire tmp7171;
  assign tmp7171 = 1'b0;
  wire tmp7172;
  assign tmp7172 = 1'b0;
  wire tmp7173;
  assign tmp7173 = (tmp7170 & tmp7171) | (tmp7170 & tmp7172) | (tmp7171 & tmp7172);
  wire tmp7174;
  assign tmp7174 = 1'b0;
  wire tmp7175;
  assign tmp7175 = 1'b0;
  wire tmp7176;
  assign tmp7176 = 1'b0;
  wire tmp7177;
  assign tmp7177 = (tmp7174 & tmp7175) | (tmp7174 & tmp7176) | (tmp7175 & tmp7176);
  wire tmp7178;
  assign tmp7178 = (tmp7169 & tmp7173) | (tmp7169 & tmp7177) | (tmp7173 & tmp7177);
  wire tmp7179;
  assign tmp7179 = 1'b0;
  wire tmp7180;
  assign tmp7180 = 1'b0;
  wire tmp7181;
  assign tmp7181 = 1'b0;
  wire tmp7182;
  assign tmp7182 = (tmp7179 & tmp7180) | (tmp7179 & tmp7181) | (tmp7180 & tmp7181);
  wire tmp7183;
  assign tmp7183 = 1'b0;
  wire tmp7184;
  assign tmp7184 = 1'b1;
  wire tmp7185;
  assign tmp7185 = 1'b0;
  wire tmp7186;
  assign tmp7186 = (tmp7183 & tmp7184) | (tmp7183 & tmp7185) | (tmp7184 & tmp7185);
  wire tmp7187;
  assign tmp7187 = 1'b0;
  wire tmp7188;
  assign tmp7188 = 1'b0;
  wire tmp7189;
  assign tmp7189 = 1'b0;
  wire tmp7190;
  assign tmp7190 = (tmp7187 & tmp7188) | (tmp7187 & tmp7189) | (tmp7188 & tmp7189);
  wire tmp7191;
  assign tmp7191 = (tmp7182 & tmp7186) | (tmp7182 & tmp7190) | (tmp7186 & tmp7190);
  wire tmp7192;
  assign tmp7192 = 1'b0;
  wire tmp7193;
  assign tmp7193 = 1'b0;
  wire tmp7194;
  assign tmp7194 = 1'b0;
  wire tmp7195;
  assign tmp7195 = (tmp7192 & tmp7193) | (tmp7192 & tmp7194) | (tmp7193 & tmp7194);
  wire tmp7196;
  assign tmp7196 = 1'b0;
  wire tmp7197;
  assign tmp7197 = 1'b0;
  wire tmp7198;
  assign tmp7198 = 1'b0;
  wire tmp7199;
  assign tmp7199 = (tmp7196 & tmp7197) | (tmp7196 & tmp7198) | (tmp7197 & tmp7198);
  wire tmp7200;
  assign tmp7200 = 1'b0;
  wire tmp7201;
  assign tmp7201 = 1'b0;
  wire tmp7202;
  assign tmp7202 = 1'b0;
  wire tmp7203;
  assign tmp7203 = (tmp7200 & tmp7201) | (tmp7200 & tmp7202) | (tmp7201 & tmp7202);
  wire tmp7204;
  assign tmp7204 = (tmp7195 & tmp7199) | (tmp7195 & tmp7203) | (tmp7199 & tmp7203);
  wire tmp7205;
  assign tmp7205 = (tmp7178 & tmp7191) | (tmp7178 & tmp7204) | (tmp7191 & tmp7204);
  wire tmp7206;
  assign tmp7206 = 1'b0;
  wire tmp7207;
  assign tmp7207 = 1'b0;
  wire tmp7208;
  assign tmp7208 = 1'b0;
  wire tmp7209;
  assign tmp7209 = (tmp7206 & tmp7207) | (tmp7206 & tmp7208) | (tmp7207 & tmp7208);
  wire tmp7210;
  assign tmp7210 = 1'b0;
  wire tmp7211;
  assign tmp7211 = 1'b1;
  wire tmp7212;
  assign tmp7212 = 1'b0;
  wire tmp7213;
  assign tmp7213 = (tmp7210 & tmp7211) | (tmp7210 & tmp7212) | (tmp7211 & tmp7212);
  wire tmp7214;
  assign tmp7214 = 1'b0;
  wire tmp7215;
  assign tmp7215 = 1'b0;
  wire tmp7216;
  assign tmp7216 = 1'b0;
  wire tmp7217;
  assign tmp7217 = (tmp7214 & tmp7215) | (tmp7214 & tmp7216) | (tmp7215 & tmp7216);
  wire tmp7218;
  assign tmp7218 = (tmp7209 & tmp7213) | (tmp7209 & tmp7217) | (tmp7213 & tmp7217);
  wire tmp7219;
  assign tmp7219 = 1'b0;
  wire tmp7220;
  assign tmp7220 = 1'b1;
  wire tmp7221;
  assign tmp7221 = 1'b0;
  wire tmp7222;
  assign tmp7222 = (tmp7219 & tmp7220) | (tmp7219 & tmp7221) | (tmp7220 & tmp7221);
  wire tmp7223;
  assign tmp7223 = 1'b1;
  wire tmp7224;
  assign tmp7224 = ~pi6;
  wire tmp7225;
  assign tmp7225 = ~pi7;
  wire tmp7226;
  assign tmp7226 = (tmp7223 & tmp7224) | (tmp7223 & tmp7225) | (tmp7224 & tmp7225);
  wire tmp7227;
  assign tmp7227 = 1'b0;
  wire tmp7228;
  assign tmp7228 = ~pi7;
  wire tmp7229;
  assign tmp7229 = 1'b0;
  wire tmp7230;
  assign tmp7230 = (tmp7227 & tmp7228) | (tmp7227 & tmp7229) | (tmp7228 & tmp7229);
  wire tmp7231;
  assign tmp7231 = (tmp7222 & tmp7226) | (tmp7222 & tmp7230) | (tmp7226 & tmp7230);
  wire tmp7232;
  assign tmp7232 = 1'b0;
  wire tmp7233;
  assign tmp7233 = 1'b0;
  wire tmp7234;
  assign tmp7234 = 1'b0;
  wire tmp7235;
  assign tmp7235 = (tmp7232 & tmp7233) | (tmp7232 & tmp7234) | (tmp7233 & tmp7234);
  wire tmp7236;
  assign tmp7236 = 1'b0;
  wire tmp7237;
  assign tmp7237 = ~pi7;
  wire tmp7238;
  assign tmp7238 = 1'b0;
  wire tmp7239;
  assign tmp7239 = (tmp7236 & tmp7237) | (tmp7236 & tmp7238) | (tmp7237 & tmp7238);
  wire tmp7240;
  assign tmp7240 = 1'b0;
  wire tmp7241;
  assign tmp7241 = 1'b0;
  wire tmp7242;
  assign tmp7242 = 1'b0;
  wire tmp7243;
  assign tmp7243 = (tmp7240 & tmp7241) | (tmp7240 & tmp7242) | (tmp7241 & tmp7242);
  wire tmp7244;
  assign tmp7244 = (tmp7235 & tmp7239) | (tmp7235 & tmp7243) | (tmp7239 & tmp7243);
  wire tmp7245;
  assign tmp7245 = (tmp7218 & tmp7231) | (tmp7218 & tmp7244) | (tmp7231 & tmp7244);
  wire tmp7246;
  assign tmp7246 = 1'b0;
  wire tmp7247;
  assign tmp7247 = 1'b0;
  wire tmp7248;
  assign tmp7248 = 1'b0;
  wire tmp7249;
  assign tmp7249 = (tmp7246 & tmp7247) | (tmp7246 & tmp7248) | (tmp7247 & tmp7248);
  wire tmp7250;
  assign tmp7250 = 1'b0;
  wire tmp7251;
  assign tmp7251 = 1'b0;
  wire tmp7252;
  assign tmp7252 = 1'b0;
  wire tmp7253;
  assign tmp7253 = (tmp7250 & tmp7251) | (tmp7250 & tmp7252) | (tmp7251 & tmp7252);
  wire tmp7254;
  assign tmp7254 = 1'b0;
  wire tmp7255;
  assign tmp7255 = 1'b0;
  wire tmp7256;
  assign tmp7256 = 1'b0;
  wire tmp7257;
  assign tmp7257 = (tmp7254 & tmp7255) | (tmp7254 & tmp7256) | (tmp7255 & tmp7256);
  wire tmp7258;
  assign tmp7258 = (tmp7249 & tmp7253) | (tmp7249 & tmp7257) | (tmp7253 & tmp7257);
  wire tmp7259;
  assign tmp7259 = 1'b0;
  wire tmp7260;
  assign tmp7260 = 1'b0;
  wire tmp7261;
  assign tmp7261 = 1'b0;
  wire tmp7262;
  assign tmp7262 = (tmp7259 & tmp7260) | (tmp7259 & tmp7261) | (tmp7260 & tmp7261);
  wire tmp7263;
  assign tmp7263 = 1'b0;
  wire tmp7264;
  assign tmp7264 = ~pi7;
  wire tmp7265;
  assign tmp7265 = 1'b0;
  wire tmp7266;
  assign tmp7266 = (tmp7263 & tmp7264) | (tmp7263 & tmp7265) | (tmp7264 & tmp7265);
  wire tmp7267;
  assign tmp7267 = 1'b0;
  wire tmp7268;
  assign tmp7268 = 1'b0;
  wire tmp7269;
  assign tmp7269 = 1'b0;
  wire tmp7270;
  assign tmp7270 = (tmp7267 & tmp7268) | (tmp7267 & tmp7269) | (tmp7268 & tmp7269);
  wire tmp7271;
  assign tmp7271 = (tmp7262 & tmp7266) | (tmp7262 & tmp7270) | (tmp7266 & tmp7270);
  wire tmp7272;
  assign tmp7272 = 1'b0;
  wire tmp7273;
  assign tmp7273 = 1'b0;
  wire tmp7274;
  assign tmp7274 = 1'b0;
  wire tmp7275;
  assign tmp7275 = (tmp7272 & tmp7273) | (tmp7272 & tmp7274) | (tmp7273 & tmp7274);
  wire tmp7276;
  assign tmp7276 = 1'b0;
  wire tmp7277;
  assign tmp7277 = 1'b0;
  wire tmp7278;
  assign tmp7278 = 1'b0;
  wire tmp7279;
  assign tmp7279 = (tmp7276 & tmp7277) | (tmp7276 & tmp7278) | (tmp7277 & tmp7278);
  wire tmp7280;
  assign tmp7280 = 1'b0;
  wire tmp7281;
  assign tmp7281 = 1'b0;
  wire tmp7282;
  assign tmp7282 = 1'b0;
  wire tmp7283;
  assign tmp7283 = (tmp7280 & tmp7281) | (tmp7280 & tmp7282) | (tmp7281 & tmp7282);
  wire tmp7284;
  assign tmp7284 = (tmp7275 & tmp7279) | (tmp7275 & tmp7283) | (tmp7279 & tmp7283);
  wire tmp7285;
  assign tmp7285 = (tmp7258 & tmp7271) | (tmp7258 & tmp7284) | (tmp7271 & tmp7284);
  wire tmp7286;
  assign tmp7286 = (tmp7205 & tmp7245) | (tmp7205 & tmp7285) | (tmp7245 & tmp7285);
  wire tmp7287;
  assign tmp7287 = (tmp7044 & tmp7165) | (tmp7044 & tmp7286) | (tmp7165 & tmp7286);
  wire tmp7288;
  assign tmp7288 = 1'b0;
  wire tmp7289;
  assign tmp7289 = 1'b0;
  wire tmp7290;
  assign tmp7290 = 1'b0;
  wire tmp7291;
  assign tmp7291 = (tmp7288 & tmp7289) | (tmp7288 & tmp7290) | (tmp7289 & tmp7290);
  wire tmp7292;
  assign tmp7292 = 1'b0;
  wire tmp7293;
  assign tmp7293 = 1'b0;
  wire tmp7294;
  assign tmp7294 = 1'b0;
  wire tmp7295;
  assign tmp7295 = (tmp7292 & tmp7293) | (tmp7292 & tmp7294) | (tmp7293 & tmp7294);
  wire tmp7296;
  assign tmp7296 = 1'b0;
  wire tmp7297;
  assign tmp7297 = 1'b0;
  wire tmp7298;
  assign tmp7298 = 1'b0;
  wire tmp7299;
  assign tmp7299 = (tmp7296 & tmp7297) | (tmp7296 & tmp7298) | (tmp7297 & tmp7298);
  wire tmp7300;
  assign tmp7300 = (tmp7291 & tmp7295) | (tmp7291 & tmp7299) | (tmp7295 & tmp7299);
  wire tmp7301;
  assign tmp7301 = 1'b0;
  wire tmp7302;
  assign tmp7302 = 1'b0;
  wire tmp7303;
  assign tmp7303 = 1'b0;
  wire tmp7304;
  assign tmp7304 = (tmp7301 & tmp7302) | (tmp7301 & tmp7303) | (tmp7302 & tmp7303);
  wire tmp7305;
  assign tmp7305 = 1'b0;
  wire tmp7306;
  assign tmp7306 = 1'b0;
  wire tmp7307;
  assign tmp7307 = 1'b0;
  wire tmp7308;
  assign tmp7308 = (tmp7305 & tmp7306) | (tmp7305 & tmp7307) | (tmp7306 & tmp7307);
  wire tmp7309;
  assign tmp7309 = 1'b0;
  wire tmp7310;
  assign tmp7310 = 1'b0;
  wire tmp7311;
  assign tmp7311 = 1'b0;
  wire tmp7312;
  assign tmp7312 = (tmp7309 & tmp7310) | (tmp7309 & tmp7311) | (tmp7310 & tmp7311);
  wire tmp7313;
  assign tmp7313 = (tmp7304 & tmp7308) | (tmp7304 & tmp7312) | (tmp7308 & tmp7312);
  wire tmp7314;
  assign tmp7314 = 1'b0;
  wire tmp7315;
  assign tmp7315 = 1'b0;
  wire tmp7316;
  assign tmp7316 = 1'b0;
  wire tmp7317;
  assign tmp7317 = (tmp7314 & tmp7315) | (tmp7314 & tmp7316) | (tmp7315 & tmp7316);
  wire tmp7318;
  assign tmp7318 = 1'b0;
  wire tmp7319;
  assign tmp7319 = 1'b0;
  wire tmp7320;
  assign tmp7320 = 1'b0;
  wire tmp7321;
  assign tmp7321 = (tmp7318 & tmp7319) | (tmp7318 & tmp7320) | (tmp7319 & tmp7320);
  wire tmp7322;
  assign tmp7322 = 1'b0;
  wire tmp7323;
  assign tmp7323 = 1'b0;
  wire tmp7324;
  assign tmp7324 = 1'b0;
  wire tmp7325;
  assign tmp7325 = (tmp7322 & tmp7323) | (tmp7322 & tmp7324) | (tmp7323 & tmp7324);
  wire tmp7326;
  assign tmp7326 = (tmp7317 & tmp7321) | (tmp7317 & tmp7325) | (tmp7321 & tmp7325);
  wire tmp7327;
  assign tmp7327 = (tmp7300 & tmp7313) | (tmp7300 & tmp7326) | (tmp7313 & tmp7326);
  wire tmp7328;
  assign tmp7328 = 1'b0;
  wire tmp7329;
  assign tmp7329 = 1'b0;
  wire tmp7330;
  assign tmp7330 = 1'b0;
  wire tmp7331;
  assign tmp7331 = (tmp7328 & tmp7329) | (tmp7328 & tmp7330) | (tmp7329 & tmp7330);
  wire tmp7332;
  assign tmp7332 = 1'b0;
  wire tmp7333;
  assign tmp7333 = 1'b0;
  wire tmp7334;
  assign tmp7334 = 1'b0;
  wire tmp7335;
  assign tmp7335 = (tmp7332 & tmp7333) | (tmp7332 & tmp7334) | (tmp7333 & tmp7334);
  wire tmp7336;
  assign tmp7336 = 1'b0;
  wire tmp7337;
  assign tmp7337 = 1'b0;
  wire tmp7338;
  assign tmp7338 = 1'b0;
  wire tmp7339;
  assign tmp7339 = (tmp7336 & tmp7337) | (tmp7336 & tmp7338) | (tmp7337 & tmp7338);
  wire tmp7340;
  assign tmp7340 = (tmp7331 & tmp7335) | (tmp7331 & tmp7339) | (tmp7335 & tmp7339);
  wire tmp7341;
  assign tmp7341 = 1'b0;
  wire tmp7342;
  assign tmp7342 = 1'b0;
  wire tmp7343;
  assign tmp7343 = 1'b0;
  wire tmp7344;
  assign tmp7344 = (tmp7341 & tmp7342) | (tmp7341 & tmp7343) | (tmp7342 & tmp7343);
  wire tmp7345;
  assign tmp7345 = 1'b0;
  wire tmp7346;
  assign tmp7346 = 1'b1;
  wire tmp7347;
  assign tmp7347 = 1'b0;
  wire tmp7348;
  assign tmp7348 = (tmp7345 & tmp7346) | (tmp7345 & tmp7347) | (tmp7346 & tmp7347);
  wire tmp7349;
  assign tmp7349 = 1'b0;
  wire tmp7350;
  assign tmp7350 = 1'b0;
  wire tmp7351;
  assign tmp7351 = 1'b0;
  wire tmp7352;
  assign tmp7352 = (tmp7349 & tmp7350) | (tmp7349 & tmp7351) | (tmp7350 & tmp7351);
  wire tmp7353;
  assign tmp7353 = (tmp7344 & tmp7348) | (tmp7344 & tmp7352) | (tmp7348 & tmp7352);
  wire tmp7354;
  assign tmp7354 = 1'b0;
  wire tmp7355;
  assign tmp7355 = 1'b0;
  wire tmp7356;
  assign tmp7356 = 1'b0;
  wire tmp7357;
  assign tmp7357 = (tmp7354 & tmp7355) | (tmp7354 & tmp7356) | (tmp7355 & tmp7356);
  wire tmp7358;
  assign tmp7358 = 1'b0;
  wire tmp7359;
  assign tmp7359 = 1'b0;
  wire tmp7360;
  assign tmp7360 = 1'b0;
  wire tmp7361;
  assign tmp7361 = (tmp7358 & tmp7359) | (tmp7358 & tmp7360) | (tmp7359 & tmp7360);
  wire tmp7362;
  assign tmp7362 = 1'b0;
  wire tmp7363;
  assign tmp7363 = 1'b0;
  wire tmp7364;
  assign tmp7364 = 1'b0;
  wire tmp7365;
  assign tmp7365 = (tmp7362 & tmp7363) | (tmp7362 & tmp7364) | (tmp7363 & tmp7364);
  wire tmp7366;
  assign tmp7366 = (tmp7357 & tmp7361) | (tmp7357 & tmp7365) | (tmp7361 & tmp7365);
  wire tmp7367;
  assign tmp7367 = (tmp7340 & tmp7353) | (tmp7340 & tmp7366) | (tmp7353 & tmp7366);
  wire tmp7368;
  assign tmp7368 = 1'b0;
  wire tmp7369;
  assign tmp7369 = 1'b0;
  wire tmp7370;
  assign tmp7370 = 1'b0;
  wire tmp7371;
  assign tmp7371 = (tmp7368 & tmp7369) | (tmp7368 & tmp7370) | (tmp7369 & tmp7370);
  wire tmp7372;
  assign tmp7372 = 1'b0;
  wire tmp7373;
  assign tmp7373 = 1'b0;
  wire tmp7374;
  assign tmp7374 = 1'b0;
  wire tmp7375;
  assign tmp7375 = (tmp7372 & tmp7373) | (tmp7372 & tmp7374) | (tmp7373 & tmp7374);
  wire tmp7376;
  assign tmp7376 = 1'b0;
  wire tmp7377;
  assign tmp7377 = 1'b0;
  wire tmp7378;
  assign tmp7378 = 1'b0;
  wire tmp7379;
  assign tmp7379 = (tmp7376 & tmp7377) | (tmp7376 & tmp7378) | (tmp7377 & tmp7378);
  wire tmp7380;
  assign tmp7380 = (tmp7371 & tmp7375) | (tmp7371 & tmp7379) | (tmp7375 & tmp7379);
  wire tmp7381;
  assign tmp7381 = 1'b0;
  wire tmp7382;
  assign tmp7382 = 1'b0;
  wire tmp7383;
  assign tmp7383 = 1'b0;
  wire tmp7384;
  assign tmp7384 = (tmp7381 & tmp7382) | (tmp7381 & tmp7383) | (tmp7382 & tmp7383);
  wire tmp7385;
  assign tmp7385 = 1'b0;
  wire tmp7386;
  assign tmp7386 = 1'b0;
  wire tmp7387;
  assign tmp7387 = 1'b0;
  wire tmp7388;
  assign tmp7388 = (tmp7385 & tmp7386) | (tmp7385 & tmp7387) | (tmp7386 & tmp7387);
  wire tmp7389;
  assign tmp7389 = 1'b0;
  wire tmp7390;
  assign tmp7390 = 1'b0;
  wire tmp7391;
  assign tmp7391 = 1'b0;
  wire tmp7392;
  assign tmp7392 = (tmp7389 & tmp7390) | (tmp7389 & tmp7391) | (tmp7390 & tmp7391);
  wire tmp7393;
  assign tmp7393 = (tmp7384 & tmp7388) | (tmp7384 & tmp7392) | (tmp7388 & tmp7392);
  wire tmp7394;
  assign tmp7394 = 1'b0;
  wire tmp7395;
  assign tmp7395 = 1'b0;
  wire tmp7396;
  assign tmp7396 = 1'b0;
  wire tmp7397;
  assign tmp7397 = (tmp7394 & tmp7395) | (tmp7394 & tmp7396) | (tmp7395 & tmp7396);
  wire tmp7398;
  assign tmp7398 = 1'b0;
  wire tmp7399;
  assign tmp7399 = 1'b0;
  wire tmp7400;
  assign tmp7400 = 1'b0;
  wire tmp7401;
  assign tmp7401 = (tmp7398 & tmp7399) | (tmp7398 & tmp7400) | (tmp7399 & tmp7400);
  wire tmp7402;
  assign tmp7402 = 1'b0;
  wire tmp7403;
  assign tmp7403 = 1'b0;
  wire tmp7404;
  assign tmp7404 = 1'b0;
  wire tmp7405;
  assign tmp7405 = (tmp7402 & tmp7403) | (tmp7402 & tmp7404) | (tmp7403 & tmp7404);
  wire tmp7406;
  assign tmp7406 = (tmp7397 & tmp7401) | (tmp7397 & tmp7405) | (tmp7401 & tmp7405);
  wire tmp7407;
  assign tmp7407 = (tmp7380 & tmp7393) | (tmp7380 & tmp7406) | (tmp7393 & tmp7406);
  wire tmp7408;
  assign tmp7408 = (tmp7327 & tmp7367) | (tmp7327 & tmp7407) | (tmp7367 & tmp7407);
  wire tmp7409;
  assign tmp7409 = 1'b0;
  wire tmp7410;
  assign tmp7410 = 1'b0;
  wire tmp7411;
  assign tmp7411 = 1'b0;
  wire tmp7412;
  assign tmp7412 = (tmp7409 & tmp7410) | (tmp7409 & tmp7411) | (tmp7410 & tmp7411);
  wire tmp7413;
  assign tmp7413 = 1'b0;
  wire tmp7414;
  assign tmp7414 = 1'b0;
  wire tmp7415;
  assign tmp7415 = 1'b0;
  wire tmp7416;
  assign tmp7416 = (tmp7413 & tmp7414) | (tmp7413 & tmp7415) | (tmp7414 & tmp7415);
  wire tmp7417;
  assign tmp7417 = 1'b0;
  wire tmp7418;
  assign tmp7418 = 1'b0;
  wire tmp7419;
  assign tmp7419 = 1'b0;
  wire tmp7420;
  assign tmp7420 = (tmp7417 & tmp7418) | (tmp7417 & tmp7419) | (tmp7418 & tmp7419);
  wire tmp7421;
  assign tmp7421 = (tmp7412 & tmp7416) | (tmp7412 & tmp7420) | (tmp7416 & tmp7420);
  wire tmp7422;
  assign tmp7422 = 1'b0;
  wire tmp7423;
  assign tmp7423 = 1'b0;
  wire tmp7424;
  assign tmp7424 = 1'b0;
  wire tmp7425;
  assign tmp7425 = (tmp7422 & tmp7423) | (tmp7422 & tmp7424) | (tmp7423 & tmp7424);
  wire tmp7426;
  assign tmp7426 = 1'b0;
  wire tmp7427;
  assign tmp7427 = 1'b1;
  wire tmp7428;
  assign tmp7428 = 1'b0;
  wire tmp7429;
  assign tmp7429 = (tmp7426 & tmp7427) | (tmp7426 & tmp7428) | (tmp7427 & tmp7428);
  wire tmp7430;
  assign tmp7430 = 1'b0;
  wire tmp7431;
  assign tmp7431 = 1'b0;
  wire tmp7432;
  assign tmp7432 = 1'b0;
  wire tmp7433;
  assign tmp7433 = (tmp7430 & tmp7431) | (tmp7430 & tmp7432) | (tmp7431 & tmp7432);
  wire tmp7434;
  assign tmp7434 = (tmp7425 & tmp7429) | (tmp7425 & tmp7433) | (tmp7429 & tmp7433);
  wire tmp7435;
  assign tmp7435 = 1'b0;
  wire tmp7436;
  assign tmp7436 = 1'b0;
  wire tmp7437;
  assign tmp7437 = 1'b0;
  wire tmp7438;
  assign tmp7438 = (tmp7435 & tmp7436) | (tmp7435 & tmp7437) | (tmp7436 & tmp7437);
  wire tmp7439;
  assign tmp7439 = 1'b0;
  wire tmp7440;
  assign tmp7440 = 1'b0;
  wire tmp7441;
  assign tmp7441 = 1'b0;
  wire tmp7442;
  assign tmp7442 = (tmp7439 & tmp7440) | (tmp7439 & tmp7441) | (tmp7440 & tmp7441);
  wire tmp7443;
  assign tmp7443 = 1'b0;
  wire tmp7444;
  assign tmp7444 = 1'b0;
  wire tmp7445;
  assign tmp7445 = 1'b0;
  wire tmp7446;
  assign tmp7446 = (tmp7443 & tmp7444) | (tmp7443 & tmp7445) | (tmp7444 & tmp7445);
  wire tmp7447;
  assign tmp7447 = (tmp7438 & tmp7442) | (tmp7438 & tmp7446) | (tmp7442 & tmp7446);
  wire tmp7448;
  assign tmp7448 = (tmp7421 & tmp7434) | (tmp7421 & tmp7447) | (tmp7434 & tmp7447);
  wire tmp7449;
  assign tmp7449 = 1'b0;
  wire tmp7450;
  assign tmp7450 = 1'b0;
  wire tmp7451;
  assign tmp7451 = 1'b0;
  wire tmp7452;
  assign tmp7452 = (tmp7449 & tmp7450) | (tmp7449 & tmp7451) | (tmp7450 & tmp7451);
  wire tmp7453;
  assign tmp7453 = 1'b0;
  wire tmp7454;
  assign tmp7454 = 1'b1;
  wire tmp7455;
  assign tmp7455 = 1'b0;
  wire tmp7456;
  assign tmp7456 = (tmp7453 & tmp7454) | (tmp7453 & tmp7455) | (tmp7454 & tmp7455);
  wire tmp7457;
  assign tmp7457 = 1'b0;
  wire tmp7458;
  assign tmp7458 = 1'b0;
  wire tmp7459;
  assign tmp7459 = 1'b0;
  wire tmp7460;
  assign tmp7460 = (tmp7457 & tmp7458) | (tmp7457 & tmp7459) | (tmp7458 & tmp7459);
  wire tmp7461;
  assign tmp7461 = (tmp7452 & tmp7456) | (tmp7452 & tmp7460) | (tmp7456 & tmp7460);
  wire tmp7462;
  assign tmp7462 = 1'b0;
  wire tmp7463;
  assign tmp7463 = 1'b1;
  wire tmp7464;
  assign tmp7464 = 1'b0;
  wire tmp7465;
  assign tmp7465 = (tmp7462 & tmp7463) | (tmp7462 & tmp7464) | (tmp7463 & tmp7464);
  wire tmp7466;
  assign tmp7466 = 1'b1;
  wire tmp7467;
  assign tmp7467 = ~pi6;
  wire tmp7468;
  assign tmp7468 = ~pi7;
  wire tmp7469;
  assign tmp7469 = (tmp7466 & tmp7467) | (tmp7466 & tmp7468) | (tmp7467 & tmp7468);
  wire tmp7470;
  assign tmp7470 = 1'b0;
  wire tmp7471;
  assign tmp7471 = ~pi7;
  wire tmp7472;
  assign tmp7472 = 1'b0;
  wire tmp7473;
  assign tmp7473 = (tmp7470 & tmp7471) | (tmp7470 & tmp7472) | (tmp7471 & tmp7472);
  wire tmp7474;
  assign tmp7474 = (tmp7465 & tmp7469) | (tmp7465 & tmp7473) | (tmp7469 & tmp7473);
  wire tmp7475;
  assign tmp7475 = 1'b0;
  wire tmp7476;
  assign tmp7476 = 1'b0;
  wire tmp7477;
  assign tmp7477 = 1'b0;
  wire tmp7478;
  assign tmp7478 = (tmp7475 & tmp7476) | (tmp7475 & tmp7477) | (tmp7476 & tmp7477);
  wire tmp7479;
  assign tmp7479 = 1'b0;
  wire tmp7480;
  assign tmp7480 = ~pi7;
  wire tmp7481;
  assign tmp7481 = 1'b0;
  wire tmp7482;
  assign tmp7482 = (tmp7479 & tmp7480) | (tmp7479 & tmp7481) | (tmp7480 & tmp7481);
  wire tmp7483;
  assign tmp7483 = 1'b0;
  wire tmp7484;
  assign tmp7484 = 1'b0;
  wire tmp7485;
  assign tmp7485 = 1'b0;
  wire tmp7486;
  assign tmp7486 = (tmp7483 & tmp7484) | (tmp7483 & tmp7485) | (tmp7484 & tmp7485);
  wire tmp7487;
  assign tmp7487 = (tmp7478 & tmp7482) | (tmp7478 & tmp7486) | (tmp7482 & tmp7486);
  wire tmp7488;
  assign tmp7488 = (tmp7461 & tmp7474) | (tmp7461 & tmp7487) | (tmp7474 & tmp7487);
  wire tmp7489;
  assign tmp7489 = 1'b0;
  wire tmp7490;
  assign tmp7490 = 1'b0;
  wire tmp7491;
  assign tmp7491 = 1'b0;
  wire tmp7492;
  assign tmp7492 = (tmp7489 & tmp7490) | (tmp7489 & tmp7491) | (tmp7490 & tmp7491);
  wire tmp7493;
  assign tmp7493 = 1'b0;
  wire tmp7494;
  assign tmp7494 = 1'b0;
  wire tmp7495;
  assign tmp7495 = 1'b0;
  wire tmp7496;
  assign tmp7496 = (tmp7493 & tmp7494) | (tmp7493 & tmp7495) | (tmp7494 & tmp7495);
  wire tmp7497;
  assign tmp7497 = 1'b0;
  wire tmp7498;
  assign tmp7498 = 1'b0;
  wire tmp7499;
  assign tmp7499 = 1'b0;
  wire tmp7500;
  assign tmp7500 = (tmp7497 & tmp7498) | (tmp7497 & tmp7499) | (tmp7498 & tmp7499);
  wire tmp7501;
  assign tmp7501 = (tmp7492 & tmp7496) | (tmp7492 & tmp7500) | (tmp7496 & tmp7500);
  wire tmp7502;
  assign tmp7502 = 1'b0;
  wire tmp7503;
  assign tmp7503 = 1'b0;
  wire tmp7504;
  assign tmp7504 = 1'b0;
  wire tmp7505;
  assign tmp7505 = (tmp7502 & tmp7503) | (tmp7502 & tmp7504) | (tmp7503 & tmp7504);
  wire tmp7506;
  assign tmp7506 = 1'b0;
  wire tmp7507;
  assign tmp7507 = ~pi7;
  wire tmp7508;
  assign tmp7508 = 1'b0;
  wire tmp7509;
  assign tmp7509 = (tmp7506 & tmp7507) | (tmp7506 & tmp7508) | (tmp7507 & tmp7508);
  wire tmp7510;
  assign tmp7510 = 1'b0;
  wire tmp7511;
  assign tmp7511 = 1'b0;
  wire tmp7512;
  assign tmp7512 = 1'b0;
  wire tmp7513;
  assign tmp7513 = (tmp7510 & tmp7511) | (tmp7510 & tmp7512) | (tmp7511 & tmp7512);
  wire tmp7514;
  assign tmp7514 = (tmp7505 & tmp7509) | (tmp7505 & tmp7513) | (tmp7509 & tmp7513);
  wire tmp7515;
  assign tmp7515 = 1'b0;
  wire tmp7516;
  assign tmp7516 = 1'b0;
  wire tmp7517;
  assign tmp7517 = 1'b0;
  wire tmp7518;
  assign tmp7518 = (tmp7515 & tmp7516) | (tmp7515 & tmp7517) | (tmp7516 & tmp7517);
  wire tmp7519;
  assign tmp7519 = 1'b0;
  wire tmp7520;
  assign tmp7520 = 1'b0;
  wire tmp7521;
  assign tmp7521 = 1'b0;
  wire tmp7522;
  assign tmp7522 = (tmp7519 & tmp7520) | (tmp7519 & tmp7521) | (tmp7520 & tmp7521);
  wire tmp7523;
  assign tmp7523 = 1'b0;
  wire tmp7524;
  assign tmp7524 = 1'b0;
  wire tmp7525;
  assign tmp7525 = 1'b0;
  wire tmp7526;
  assign tmp7526 = (tmp7523 & tmp7524) | (tmp7523 & tmp7525) | (tmp7524 & tmp7525);
  wire tmp7527;
  assign tmp7527 = (tmp7518 & tmp7522) | (tmp7518 & tmp7526) | (tmp7522 & tmp7526);
  wire tmp7528;
  assign tmp7528 = (tmp7501 & tmp7514) | (tmp7501 & tmp7527) | (tmp7514 & tmp7527);
  wire tmp7529;
  assign tmp7529 = (tmp7448 & tmp7488) | (tmp7448 & tmp7528) | (tmp7488 & tmp7528);
  wire tmp7530;
  assign tmp7530 = 1'b0;
  wire tmp7531;
  assign tmp7531 = 1'b0;
  wire tmp7532;
  assign tmp7532 = 1'b0;
  wire tmp7533;
  assign tmp7533 = (tmp7530 & tmp7531) | (tmp7530 & tmp7532) | (tmp7531 & tmp7532);
  wire tmp7534;
  assign tmp7534 = 1'b0;
  wire tmp7535;
  assign tmp7535 = 1'b0;
  wire tmp7536;
  assign tmp7536 = 1'b0;
  wire tmp7537;
  assign tmp7537 = (tmp7534 & tmp7535) | (tmp7534 & tmp7536) | (tmp7535 & tmp7536);
  wire tmp7538;
  assign tmp7538 = 1'b0;
  wire tmp7539;
  assign tmp7539 = 1'b0;
  wire tmp7540;
  assign tmp7540 = 1'b0;
  wire tmp7541;
  assign tmp7541 = (tmp7538 & tmp7539) | (tmp7538 & tmp7540) | (tmp7539 & tmp7540);
  wire tmp7542;
  assign tmp7542 = (tmp7533 & tmp7537) | (tmp7533 & tmp7541) | (tmp7537 & tmp7541);
  wire tmp7543;
  assign tmp7543 = 1'b0;
  wire tmp7544;
  assign tmp7544 = 1'b0;
  wire tmp7545;
  assign tmp7545 = 1'b0;
  wire tmp7546;
  assign tmp7546 = (tmp7543 & tmp7544) | (tmp7543 & tmp7545) | (tmp7544 & tmp7545);
  wire tmp7547;
  assign tmp7547 = 1'b0;
  wire tmp7548;
  assign tmp7548 = 1'b0;
  wire tmp7549;
  assign tmp7549 = 1'b0;
  wire tmp7550;
  assign tmp7550 = (tmp7547 & tmp7548) | (tmp7547 & tmp7549) | (tmp7548 & tmp7549);
  wire tmp7551;
  assign tmp7551 = 1'b0;
  wire tmp7552;
  assign tmp7552 = 1'b0;
  wire tmp7553;
  assign tmp7553 = 1'b0;
  wire tmp7554;
  assign tmp7554 = (tmp7551 & tmp7552) | (tmp7551 & tmp7553) | (tmp7552 & tmp7553);
  wire tmp7555;
  assign tmp7555 = (tmp7546 & tmp7550) | (tmp7546 & tmp7554) | (tmp7550 & tmp7554);
  wire tmp7556;
  assign tmp7556 = 1'b0;
  wire tmp7557;
  assign tmp7557 = 1'b0;
  wire tmp7558;
  assign tmp7558 = 1'b0;
  wire tmp7559;
  assign tmp7559 = (tmp7556 & tmp7557) | (tmp7556 & tmp7558) | (tmp7557 & tmp7558);
  wire tmp7560;
  assign tmp7560 = 1'b0;
  wire tmp7561;
  assign tmp7561 = 1'b0;
  wire tmp7562;
  assign tmp7562 = 1'b0;
  wire tmp7563;
  assign tmp7563 = (tmp7560 & tmp7561) | (tmp7560 & tmp7562) | (tmp7561 & tmp7562);
  wire tmp7564;
  assign tmp7564 = 1'b0;
  wire tmp7565;
  assign tmp7565 = 1'b0;
  wire tmp7566;
  assign tmp7566 = 1'b0;
  wire tmp7567;
  assign tmp7567 = (tmp7564 & tmp7565) | (tmp7564 & tmp7566) | (tmp7565 & tmp7566);
  wire tmp7568;
  assign tmp7568 = (tmp7559 & tmp7563) | (tmp7559 & tmp7567) | (tmp7563 & tmp7567);
  wire tmp7569;
  assign tmp7569 = (tmp7542 & tmp7555) | (tmp7542 & tmp7568) | (tmp7555 & tmp7568);
  wire tmp7570;
  assign tmp7570 = 1'b0;
  wire tmp7571;
  assign tmp7571 = 1'b0;
  wire tmp7572;
  assign tmp7572 = 1'b0;
  wire tmp7573;
  assign tmp7573 = (tmp7570 & tmp7571) | (tmp7570 & tmp7572) | (tmp7571 & tmp7572);
  wire tmp7574;
  assign tmp7574 = 1'b0;
  wire tmp7575;
  assign tmp7575 = 1'b0;
  wire tmp7576;
  assign tmp7576 = 1'b0;
  wire tmp7577;
  assign tmp7577 = (tmp7574 & tmp7575) | (tmp7574 & tmp7576) | (tmp7575 & tmp7576);
  wire tmp7578;
  assign tmp7578 = 1'b0;
  wire tmp7579;
  assign tmp7579 = 1'b0;
  wire tmp7580;
  assign tmp7580 = 1'b0;
  wire tmp7581;
  assign tmp7581 = (tmp7578 & tmp7579) | (tmp7578 & tmp7580) | (tmp7579 & tmp7580);
  wire tmp7582;
  assign tmp7582 = (tmp7573 & tmp7577) | (tmp7573 & tmp7581) | (tmp7577 & tmp7581);
  wire tmp7583;
  assign tmp7583 = 1'b0;
  wire tmp7584;
  assign tmp7584 = 1'b0;
  wire tmp7585;
  assign tmp7585 = 1'b0;
  wire tmp7586;
  assign tmp7586 = (tmp7583 & tmp7584) | (tmp7583 & tmp7585) | (tmp7584 & tmp7585);
  wire tmp7587;
  assign tmp7587 = 1'b0;
  wire tmp7588;
  assign tmp7588 = ~pi7;
  wire tmp7589;
  assign tmp7589 = 1'b0;
  wire tmp7590;
  assign tmp7590 = (tmp7587 & tmp7588) | (tmp7587 & tmp7589) | (tmp7588 & tmp7589);
  wire tmp7591;
  assign tmp7591 = 1'b0;
  wire tmp7592;
  assign tmp7592 = 1'b0;
  wire tmp7593;
  assign tmp7593 = 1'b0;
  wire tmp7594;
  assign tmp7594 = (tmp7591 & tmp7592) | (tmp7591 & tmp7593) | (tmp7592 & tmp7593);
  wire tmp7595;
  assign tmp7595 = (tmp7586 & tmp7590) | (tmp7586 & tmp7594) | (tmp7590 & tmp7594);
  wire tmp7596;
  assign tmp7596 = 1'b0;
  wire tmp7597;
  assign tmp7597 = 1'b0;
  wire tmp7598;
  assign tmp7598 = 1'b0;
  wire tmp7599;
  assign tmp7599 = (tmp7596 & tmp7597) | (tmp7596 & tmp7598) | (tmp7597 & tmp7598);
  wire tmp7600;
  assign tmp7600 = 1'b0;
  wire tmp7601;
  assign tmp7601 = 1'b0;
  wire tmp7602;
  assign tmp7602 = 1'b0;
  wire tmp7603;
  assign tmp7603 = (tmp7600 & tmp7601) | (tmp7600 & tmp7602) | (tmp7601 & tmp7602);
  wire tmp7604;
  assign tmp7604 = 1'b0;
  wire tmp7605;
  assign tmp7605 = 1'b0;
  wire tmp7606;
  assign tmp7606 = 1'b0;
  wire tmp7607;
  assign tmp7607 = (tmp7604 & tmp7605) | (tmp7604 & tmp7606) | (tmp7605 & tmp7606);
  wire tmp7608;
  assign tmp7608 = (tmp7599 & tmp7603) | (tmp7599 & tmp7607) | (tmp7603 & tmp7607);
  wire tmp7609;
  assign tmp7609 = (tmp7582 & tmp7595) | (tmp7582 & tmp7608) | (tmp7595 & tmp7608);
  wire tmp7610;
  assign tmp7610 = 1'b0;
  wire tmp7611;
  assign tmp7611 = 1'b0;
  wire tmp7612;
  assign tmp7612 = 1'b0;
  wire tmp7613;
  assign tmp7613 = (tmp7610 & tmp7611) | (tmp7610 & tmp7612) | (tmp7611 & tmp7612);
  wire tmp7614;
  assign tmp7614 = 1'b0;
  wire tmp7615;
  assign tmp7615 = 1'b0;
  wire tmp7616;
  assign tmp7616 = 1'b0;
  wire tmp7617;
  assign tmp7617 = (tmp7614 & tmp7615) | (tmp7614 & tmp7616) | (tmp7615 & tmp7616);
  wire tmp7618;
  assign tmp7618 = 1'b0;
  wire tmp7619;
  assign tmp7619 = 1'b0;
  wire tmp7620;
  assign tmp7620 = 1'b0;
  wire tmp7621;
  assign tmp7621 = (tmp7618 & tmp7619) | (tmp7618 & tmp7620) | (tmp7619 & tmp7620);
  wire tmp7622;
  assign tmp7622 = (tmp7613 & tmp7617) | (tmp7613 & tmp7621) | (tmp7617 & tmp7621);
  wire tmp7623;
  assign tmp7623 = 1'b0;
  wire tmp7624;
  assign tmp7624 = 1'b0;
  wire tmp7625;
  assign tmp7625 = 1'b0;
  wire tmp7626;
  assign tmp7626 = (tmp7623 & tmp7624) | (tmp7623 & tmp7625) | (tmp7624 & tmp7625);
  wire tmp7627;
  assign tmp7627 = 1'b0;
  wire tmp7628;
  assign tmp7628 = 1'b0;
  wire tmp7629;
  assign tmp7629 = 1'b0;
  wire tmp7630;
  assign tmp7630 = (tmp7627 & tmp7628) | (tmp7627 & tmp7629) | (tmp7628 & tmp7629);
  wire tmp7631;
  assign tmp7631 = 1'b0;
  wire tmp7632;
  assign tmp7632 = 1'b0;
  wire tmp7633;
  assign tmp7633 = 1'b0;
  wire tmp7634;
  assign tmp7634 = (tmp7631 & tmp7632) | (tmp7631 & tmp7633) | (tmp7632 & tmp7633);
  wire tmp7635;
  assign tmp7635 = (tmp7626 & tmp7630) | (tmp7626 & tmp7634) | (tmp7630 & tmp7634);
  wire tmp7636;
  assign tmp7636 = 1'b0;
  wire tmp7637;
  assign tmp7637 = 1'b0;
  wire tmp7638;
  assign tmp7638 = 1'b0;
  wire tmp7639;
  assign tmp7639 = (tmp7636 & tmp7637) | (tmp7636 & tmp7638) | (tmp7637 & tmp7638);
  wire tmp7640;
  assign tmp7640 = 1'b0;
  wire tmp7641;
  assign tmp7641 = 1'b0;
  wire tmp7642;
  assign tmp7642 = 1'b0;
  wire tmp7643;
  assign tmp7643 = (tmp7640 & tmp7641) | (tmp7640 & tmp7642) | (tmp7641 & tmp7642);
  wire tmp7644;
  assign tmp7644 = 1'b0;
  wire tmp7645;
  assign tmp7645 = 1'b0;
  wire tmp7646;
  assign tmp7646 = 1'b0;
  wire tmp7647;
  assign tmp7647 = (tmp7644 & tmp7645) | (tmp7644 & tmp7646) | (tmp7645 & tmp7646);
  wire tmp7648;
  assign tmp7648 = (tmp7639 & tmp7643) | (tmp7639 & tmp7647) | (tmp7643 & tmp7647);
  wire tmp7649;
  assign tmp7649 = (tmp7622 & tmp7635) | (tmp7622 & tmp7648) | (tmp7635 & tmp7648);
  wire tmp7650;
  assign tmp7650 = (tmp7569 & tmp7609) | (tmp7569 & tmp7649) | (tmp7609 & tmp7649);
  wire tmp7651;
  assign tmp7651 = (tmp7408 & tmp7529) | (tmp7408 & tmp7650) | (tmp7529 & tmp7650);
  wire tmp7652;
  assign tmp7652 = (tmp6923 & tmp7287) | (tmp6923 & tmp7651) | (tmp7287 & tmp7651);
  wire tmp7653;
  assign tmp7653 = 1'b0;
  wire tmp7654;
  assign tmp7654 = 1'b0;
  wire tmp7655;
  assign tmp7655 = 1'b0;
  wire tmp7656;
  assign tmp7656 = (tmp7653 & tmp7654) | (tmp7653 & tmp7655) | (tmp7654 & tmp7655);
  wire tmp7657;
  assign tmp7657 = 1'b0;
  wire tmp7658;
  assign tmp7658 = 1'b0;
  wire tmp7659;
  assign tmp7659 = 1'b0;
  wire tmp7660;
  assign tmp7660 = (tmp7657 & tmp7658) | (tmp7657 & tmp7659) | (tmp7658 & tmp7659);
  wire tmp7661;
  assign tmp7661 = 1'b0;
  wire tmp7662;
  assign tmp7662 = 1'b0;
  wire tmp7663;
  assign tmp7663 = 1'b0;
  wire tmp7664;
  assign tmp7664 = (tmp7661 & tmp7662) | (tmp7661 & tmp7663) | (tmp7662 & tmp7663);
  wire tmp7665;
  assign tmp7665 = (tmp7656 & tmp7660) | (tmp7656 & tmp7664) | (tmp7660 & tmp7664);
  wire tmp7666;
  assign tmp7666 = 1'b0;
  wire tmp7667;
  assign tmp7667 = 1'b0;
  wire tmp7668;
  assign tmp7668 = 1'b0;
  wire tmp7669;
  assign tmp7669 = (tmp7666 & tmp7667) | (tmp7666 & tmp7668) | (tmp7667 & tmp7668);
  wire tmp7670;
  assign tmp7670 = 1'b0;
  wire tmp7671;
  assign tmp7671 = 1'b1;
  wire tmp7672;
  assign tmp7672 = 1'b0;
  wire tmp7673;
  assign tmp7673 = (tmp7670 & tmp7671) | (tmp7670 & tmp7672) | (tmp7671 & tmp7672);
  wire tmp7674;
  assign tmp7674 = 1'b0;
  wire tmp7675;
  assign tmp7675 = 1'b0;
  wire tmp7676;
  assign tmp7676 = 1'b0;
  wire tmp7677;
  assign tmp7677 = (tmp7674 & tmp7675) | (tmp7674 & tmp7676) | (tmp7675 & tmp7676);
  wire tmp7678;
  assign tmp7678 = (tmp7669 & tmp7673) | (tmp7669 & tmp7677) | (tmp7673 & tmp7677);
  wire tmp7679;
  assign tmp7679 = 1'b0;
  wire tmp7680;
  assign tmp7680 = 1'b0;
  wire tmp7681;
  assign tmp7681 = 1'b0;
  wire tmp7682;
  assign tmp7682 = (tmp7679 & tmp7680) | (tmp7679 & tmp7681) | (tmp7680 & tmp7681);
  wire tmp7683;
  assign tmp7683 = 1'b0;
  wire tmp7684;
  assign tmp7684 = 1'b0;
  wire tmp7685;
  assign tmp7685 = 1'b0;
  wire tmp7686;
  assign tmp7686 = (tmp7683 & tmp7684) | (tmp7683 & tmp7685) | (tmp7684 & tmp7685);
  wire tmp7687;
  assign tmp7687 = 1'b0;
  wire tmp7688;
  assign tmp7688 = 1'b0;
  wire tmp7689;
  assign tmp7689 = 1'b0;
  wire tmp7690;
  assign tmp7690 = (tmp7687 & tmp7688) | (tmp7687 & tmp7689) | (tmp7688 & tmp7689);
  wire tmp7691;
  assign tmp7691 = (tmp7682 & tmp7686) | (tmp7682 & tmp7690) | (tmp7686 & tmp7690);
  wire tmp7692;
  assign tmp7692 = (tmp7665 & tmp7678) | (tmp7665 & tmp7691) | (tmp7678 & tmp7691);
  wire tmp7693;
  assign tmp7693 = 1'b0;
  wire tmp7694;
  assign tmp7694 = 1'b0;
  wire tmp7695;
  assign tmp7695 = 1'b0;
  wire tmp7696;
  assign tmp7696 = (tmp7693 & tmp7694) | (tmp7693 & tmp7695) | (tmp7694 & tmp7695);
  wire tmp7697;
  assign tmp7697 = 1'b0;
  wire tmp7698;
  assign tmp7698 = 1'b1;
  wire tmp7699;
  assign tmp7699 = 1'b0;
  wire tmp7700;
  assign tmp7700 = (tmp7697 & tmp7698) | (tmp7697 & tmp7699) | (tmp7698 & tmp7699);
  wire tmp7701;
  assign tmp7701 = 1'b0;
  wire tmp7702;
  assign tmp7702 = 1'b0;
  wire tmp7703;
  assign tmp7703 = 1'b0;
  wire tmp7704;
  assign tmp7704 = (tmp7701 & tmp7702) | (tmp7701 & tmp7703) | (tmp7702 & tmp7703);
  wire tmp7705;
  assign tmp7705 = (tmp7696 & tmp7700) | (tmp7696 & tmp7704) | (tmp7700 & tmp7704);
  wire tmp7706;
  assign tmp7706 = 1'b0;
  wire tmp7707;
  assign tmp7707 = 1'b1;
  wire tmp7708;
  assign tmp7708 = 1'b0;
  wire tmp7709;
  assign tmp7709 = (tmp7706 & tmp7707) | (tmp7706 & tmp7708) | (tmp7707 & tmp7708);
  wire tmp7710;
  assign tmp7710 = 1'b1;
  wire tmp7711;
  assign tmp7711 = 1'b1;
  wire tmp7712;
  assign tmp7712 = 1'b1;
  wire tmp7713;
  assign tmp7713 = (tmp7710 & tmp7711) | (tmp7710 & tmp7712) | (tmp7711 & tmp7712);
  wire tmp7714;
  assign tmp7714 = 1'b0;
  wire tmp7715;
  assign tmp7715 = 1'b1;
  wire tmp7716;
  assign tmp7716 = 1'b0;
  wire tmp7717;
  assign tmp7717 = (tmp7714 & tmp7715) | (tmp7714 & tmp7716) | (tmp7715 & tmp7716);
  wire tmp7718;
  assign tmp7718 = (tmp7709 & tmp7713) | (tmp7709 & tmp7717) | (tmp7713 & tmp7717);
  wire tmp7719;
  assign tmp7719 = 1'b0;
  wire tmp7720;
  assign tmp7720 = 1'b0;
  wire tmp7721;
  assign tmp7721 = 1'b0;
  wire tmp7722;
  assign tmp7722 = (tmp7719 & tmp7720) | (tmp7719 & tmp7721) | (tmp7720 & tmp7721);
  wire tmp7723;
  assign tmp7723 = 1'b0;
  wire tmp7724;
  assign tmp7724 = 1'b1;
  wire tmp7725;
  assign tmp7725 = 1'b0;
  wire tmp7726;
  assign tmp7726 = (tmp7723 & tmp7724) | (tmp7723 & tmp7725) | (tmp7724 & tmp7725);
  wire tmp7727;
  assign tmp7727 = 1'b0;
  wire tmp7728;
  assign tmp7728 = 1'b0;
  wire tmp7729;
  assign tmp7729 = 1'b0;
  wire tmp7730;
  assign tmp7730 = (tmp7727 & tmp7728) | (tmp7727 & tmp7729) | (tmp7728 & tmp7729);
  wire tmp7731;
  assign tmp7731 = (tmp7722 & tmp7726) | (tmp7722 & tmp7730) | (tmp7726 & tmp7730);
  wire tmp7732;
  assign tmp7732 = (tmp7705 & tmp7718) | (tmp7705 & tmp7731) | (tmp7718 & tmp7731);
  wire tmp7733;
  assign tmp7733 = 1'b0;
  wire tmp7734;
  assign tmp7734 = 1'b0;
  wire tmp7735;
  assign tmp7735 = 1'b0;
  wire tmp7736;
  assign tmp7736 = (tmp7733 & tmp7734) | (tmp7733 & tmp7735) | (tmp7734 & tmp7735);
  wire tmp7737;
  assign tmp7737 = 1'b0;
  wire tmp7738;
  assign tmp7738 = 1'b0;
  wire tmp7739;
  assign tmp7739 = 1'b0;
  wire tmp7740;
  assign tmp7740 = (tmp7737 & tmp7738) | (tmp7737 & tmp7739) | (tmp7738 & tmp7739);
  wire tmp7741;
  assign tmp7741 = 1'b0;
  wire tmp7742;
  assign tmp7742 = 1'b0;
  wire tmp7743;
  assign tmp7743 = 1'b0;
  wire tmp7744;
  assign tmp7744 = (tmp7741 & tmp7742) | (tmp7741 & tmp7743) | (tmp7742 & tmp7743);
  wire tmp7745;
  assign tmp7745 = (tmp7736 & tmp7740) | (tmp7736 & tmp7744) | (tmp7740 & tmp7744);
  wire tmp7746;
  assign tmp7746 = 1'b0;
  wire tmp7747;
  assign tmp7747 = 1'b0;
  wire tmp7748;
  assign tmp7748 = 1'b0;
  wire tmp7749;
  assign tmp7749 = (tmp7746 & tmp7747) | (tmp7746 & tmp7748) | (tmp7747 & tmp7748);
  wire tmp7750;
  assign tmp7750 = 1'b0;
  wire tmp7751;
  assign tmp7751 = 1'b1;
  wire tmp7752;
  assign tmp7752 = 1'b0;
  wire tmp7753;
  assign tmp7753 = (tmp7750 & tmp7751) | (tmp7750 & tmp7752) | (tmp7751 & tmp7752);
  wire tmp7754;
  assign tmp7754 = 1'b0;
  wire tmp7755;
  assign tmp7755 = 1'b0;
  wire tmp7756;
  assign tmp7756 = 1'b0;
  wire tmp7757;
  assign tmp7757 = (tmp7754 & tmp7755) | (tmp7754 & tmp7756) | (tmp7755 & tmp7756);
  wire tmp7758;
  assign tmp7758 = (tmp7749 & tmp7753) | (tmp7749 & tmp7757) | (tmp7753 & tmp7757);
  wire tmp7759;
  assign tmp7759 = 1'b0;
  wire tmp7760;
  assign tmp7760 = 1'b0;
  wire tmp7761;
  assign tmp7761 = 1'b0;
  wire tmp7762;
  assign tmp7762 = (tmp7759 & tmp7760) | (tmp7759 & tmp7761) | (tmp7760 & tmp7761);
  wire tmp7763;
  assign tmp7763 = 1'b0;
  wire tmp7764;
  assign tmp7764 = 1'b0;
  wire tmp7765;
  assign tmp7765 = 1'b0;
  wire tmp7766;
  assign tmp7766 = (tmp7763 & tmp7764) | (tmp7763 & tmp7765) | (tmp7764 & tmp7765);
  wire tmp7767;
  assign tmp7767 = 1'b0;
  wire tmp7768;
  assign tmp7768 = 1'b0;
  wire tmp7769;
  assign tmp7769 = 1'b0;
  wire tmp7770;
  assign tmp7770 = (tmp7767 & tmp7768) | (tmp7767 & tmp7769) | (tmp7768 & tmp7769);
  wire tmp7771;
  assign tmp7771 = (tmp7762 & tmp7766) | (tmp7762 & tmp7770) | (tmp7766 & tmp7770);
  wire tmp7772;
  assign tmp7772 = (tmp7745 & tmp7758) | (tmp7745 & tmp7771) | (tmp7758 & tmp7771);
  wire tmp7773;
  assign tmp7773 = (tmp7692 & tmp7732) | (tmp7692 & tmp7772) | (tmp7732 & tmp7772);
  wire tmp7774;
  assign tmp7774 = 1'b0;
  wire tmp7775;
  assign tmp7775 = 1'b0;
  wire tmp7776;
  assign tmp7776 = 1'b0;
  wire tmp7777;
  assign tmp7777 = (tmp7774 & tmp7775) | (tmp7774 & tmp7776) | (tmp7775 & tmp7776);
  wire tmp7778;
  assign tmp7778 = 1'b0;
  wire tmp7779;
  assign tmp7779 = 1'b1;
  wire tmp7780;
  assign tmp7780 = 1'b0;
  wire tmp7781;
  assign tmp7781 = (tmp7778 & tmp7779) | (tmp7778 & tmp7780) | (tmp7779 & tmp7780);
  wire tmp7782;
  assign tmp7782 = 1'b0;
  wire tmp7783;
  assign tmp7783 = 1'b0;
  wire tmp7784;
  assign tmp7784 = 1'b0;
  wire tmp7785;
  assign tmp7785 = (tmp7782 & tmp7783) | (tmp7782 & tmp7784) | (tmp7783 & tmp7784);
  wire tmp7786;
  assign tmp7786 = (tmp7777 & tmp7781) | (tmp7777 & tmp7785) | (tmp7781 & tmp7785);
  wire tmp7787;
  assign tmp7787 = 1'b0;
  wire tmp7788;
  assign tmp7788 = 1'b1;
  wire tmp7789;
  assign tmp7789 = 1'b0;
  wire tmp7790;
  assign tmp7790 = (tmp7787 & tmp7788) | (tmp7787 & tmp7789) | (tmp7788 & tmp7789);
  wire tmp7791;
  assign tmp7791 = 1'b1;
  wire tmp7792;
  assign tmp7792 = 1'b1;
  wire tmp7793;
  assign tmp7793 = 1'b1;
  wire tmp7794;
  assign tmp7794 = (tmp7791 & tmp7792) | (tmp7791 & tmp7793) | (tmp7792 & tmp7793);
  wire tmp7795;
  assign tmp7795 = 1'b0;
  wire tmp7796;
  assign tmp7796 = 1'b1;
  wire tmp7797;
  assign tmp7797 = 1'b0;
  wire tmp7798;
  assign tmp7798 = (tmp7795 & tmp7796) | (tmp7795 & tmp7797) | (tmp7796 & tmp7797);
  wire tmp7799;
  assign tmp7799 = (tmp7790 & tmp7794) | (tmp7790 & tmp7798) | (tmp7794 & tmp7798);
  wire tmp7800;
  assign tmp7800 = 1'b0;
  wire tmp7801;
  assign tmp7801 = 1'b0;
  wire tmp7802;
  assign tmp7802 = 1'b0;
  wire tmp7803;
  assign tmp7803 = (tmp7800 & tmp7801) | (tmp7800 & tmp7802) | (tmp7801 & tmp7802);
  wire tmp7804;
  assign tmp7804 = 1'b0;
  wire tmp7805;
  assign tmp7805 = 1'b1;
  wire tmp7806;
  assign tmp7806 = 1'b0;
  wire tmp7807;
  assign tmp7807 = (tmp7804 & tmp7805) | (tmp7804 & tmp7806) | (tmp7805 & tmp7806);
  wire tmp7808;
  assign tmp7808 = 1'b0;
  wire tmp7809;
  assign tmp7809 = 1'b0;
  wire tmp7810;
  assign tmp7810 = 1'b0;
  wire tmp7811;
  assign tmp7811 = (tmp7808 & tmp7809) | (tmp7808 & tmp7810) | (tmp7809 & tmp7810);
  wire tmp7812;
  assign tmp7812 = (tmp7803 & tmp7807) | (tmp7803 & tmp7811) | (tmp7807 & tmp7811);
  wire tmp7813;
  assign tmp7813 = (tmp7786 & tmp7799) | (tmp7786 & tmp7812) | (tmp7799 & tmp7812);
  wire tmp7814;
  assign tmp7814 = 1'b0;
  wire tmp7815;
  assign tmp7815 = 1'b1;
  wire tmp7816;
  assign tmp7816 = 1'b0;
  wire tmp7817;
  assign tmp7817 = (tmp7814 & tmp7815) | (tmp7814 & tmp7816) | (tmp7815 & tmp7816);
  wire tmp7818;
  assign tmp7818 = 1'b1;
  wire tmp7819;
  assign tmp7819 = 1'b1;
  wire tmp7820;
  assign tmp7820 = 1'b1;
  wire tmp7821;
  assign tmp7821 = (tmp7818 & tmp7819) | (tmp7818 & tmp7820) | (tmp7819 & tmp7820);
  wire tmp7822;
  assign tmp7822 = 1'b0;
  wire tmp7823;
  assign tmp7823 = 1'b1;
  wire tmp7824;
  assign tmp7824 = 1'b0;
  wire tmp7825;
  assign tmp7825 = (tmp7822 & tmp7823) | (tmp7822 & tmp7824) | (tmp7823 & tmp7824);
  wire tmp7826;
  assign tmp7826 = (tmp7817 & tmp7821) | (tmp7817 & tmp7825) | (tmp7821 & tmp7825);
  wire tmp7827;
  assign tmp7827 = 1'b1;
  wire tmp7828;
  assign tmp7828 = 1'b1;
  wire tmp7829;
  assign tmp7829 = 1'b1;
  wire tmp7830;
  assign tmp7830 = (tmp7827 & tmp7828) | (tmp7827 & tmp7829) | (tmp7828 & tmp7829);
  wire tmp7831;
  assign tmp7831 = 1'b1;
  wire tmp7832;
  assign tmp7832 = ~pi5;
  wire tmp7833;
  assign tmp7833 = ~pi6;
  wire tmp7834;
  assign tmp7834 = (tmp7831 & tmp7832) | (tmp7831 & tmp7833) | (tmp7832 & tmp7833);
  wire tmp7835;
  assign tmp7835 = 1'b1;
  wire tmp7836;
  assign tmp7836 = ~pi6;
  wire tmp7837;
  assign tmp7837 = ~pi7;
  wire tmp7838;
  assign tmp7838 = (tmp7835 & tmp7836) | (tmp7835 & tmp7837) | (tmp7836 & tmp7837);
  wire tmp7839;
  assign tmp7839 = (tmp7830 & tmp7834) | (tmp7830 & tmp7838) | (tmp7834 & tmp7838);
  wire tmp7840;
  assign tmp7840 = 1'b0;
  wire tmp7841;
  assign tmp7841 = 1'b1;
  wire tmp7842;
  assign tmp7842 = 1'b0;
  wire tmp7843;
  assign tmp7843 = (tmp7840 & tmp7841) | (tmp7840 & tmp7842) | (tmp7841 & tmp7842);
  wire tmp7844;
  assign tmp7844 = 1'b1;
  wire tmp7845;
  assign tmp7845 = ~pi6;
  wire tmp7846;
  assign tmp7846 = ~pi7;
  wire tmp7847;
  assign tmp7847 = (tmp7844 & tmp7845) | (tmp7844 & tmp7846) | (tmp7845 & tmp7846);
  wire tmp7848;
  assign tmp7848 = 1'b0;
  wire tmp7849;
  assign tmp7849 = ~pi7;
  wire tmp7850;
  assign tmp7850 = 1'b0;
  wire tmp7851;
  assign tmp7851 = (tmp7848 & tmp7849) | (tmp7848 & tmp7850) | (tmp7849 & tmp7850);
  wire tmp7852;
  assign tmp7852 = (tmp7843 & tmp7847) | (tmp7843 & tmp7851) | (tmp7847 & tmp7851);
  wire tmp7853;
  assign tmp7853 = (tmp7826 & tmp7839) | (tmp7826 & tmp7852) | (tmp7839 & tmp7852);
  wire tmp7854;
  assign tmp7854 = 1'b0;
  wire tmp7855;
  assign tmp7855 = 1'b0;
  wire tmp7856;
  assign tmp7856 = 1'b0;
  wire tmp7857;
  assign tmp7857 = (tmp7854 & tmp7855) | (tmp7854 & tmp7856) | (tmp7855 & tmp7856);
  wire tmp7858;
  assign tmp7858 = 1'b0;
  wire tmp7859;
  assign tmp7859 = 1'b1;
  wire tmp7860;
  assign tmp7860 = 1'b0;
  wire tmp7861;
  assign tmp7861 = (tmp7858 & tmp7859) | (tmp7858 & tmp7860) | (tmp7859 & tmp7860);
  wire tmp7862;
  assign tmp7862 = 1'b0;
  wire tmp7863;
  assign tmp7863 = 1'b0;
  wire tmp7864;
  assign tmp7864 = 1'b0;
  wire tmp7865;
  assign tmp7865 = (tmp7862 & tmp7863) | (tmp7862 & tmp7864) | (tmp7863 & tmp7864);
  wire tmp7866;
  assign tmp7866 = (tmp7857 & tmp7861) | (tmp7857 & tmp7865) | (tmp7861 & tmp7865);
  wire tmp7867;
  assign tmp7867 = 1'b0;
  wire tmp7868;
  assign tmp7868 = 1'b1;
  wire tmp7869;
  assign tmp7869 = 1'b0;
  wire tmp7870;
  assign tmp7870 = (tmp7867 & tmp7868) | (tmp7867 & tmp7869) | (tmp7868 & tmp7869);
  wire tmp7871;
  assign tmp7871 = 1'b1;
  wire tmp7872;
  assign tmp7872 = ~pi6;
  wire tmp7873;
  assign tmp7873 = ~pi7;
  wire tmp7874;
  assign tmp7874 = (tmp7871 & tmp7872) | (tmp7871 & tmp7873) | (tmp7872 & tmp7873);
  wire tmp7875;
  assign tmp7875 = 1'b0;
  wire tmp7876;
  assign tmp7876 = ~pi7;
  wire tmp7877;
  assign tmp7877 = 1'b0;
  wire tmp7878;
  assign tmp7878 = (tmp7875 & tmp7876) | (tmp7875 & tmp7877) | (tmp7876 & tmp7877);
  wire tmp7879;
  assign tmp7879 = (tmp7870 & tmp7874) | (tmp7870 & tmp7878) | (tmp7874 & tmp7878);
  wire tmp7880;
  assign tmp7880 = 1'b0;
  wire tmp7881;
  assign tmp7881 = 1'b0;
  wire tmp7882;
  assign tmp7882 = 1'b0;
  wire tmp7883;
  assign tmp7883 = (tmp7880 & tmp7881) | (tmp7880 & tmp7882) | (tmp7881 & tmp7882);
  wire tmp7884;
  assign tmp7884 = 1'b0;
  wire tmp7885;
  assign tmp7885 = ~pi7;
  wire tmp7886;
  assign tmp7886 = 1'b0;
  wire tmp7887;
  assign tmp7887 = (tmp7884 & tmp7885) | (tmp7884 & tmp7886) | (tmp7885 & tmp7886);
  wire tmp7888;
  assign tmp7888 = 1'b0;
  wire tmp7889;
  assign tmp7889 = 1'b0;
  wire tmp7890;
  assign tmp7890 = 1'b0;
  wire tmp7891;
  assign tmp7891 = (tmp7888 & tmp7889) | (tmp7888 & tmp7890) | (tmp7889 & tmp7890);
  wire tmp7892;
  assign tmp7892 = (tmp7883 & tmp7887) | (tmp7883 & tmp7891) | (tmp7887 & tmp7891);
  wire tmp7893;
  assign tmp7893 = (tmp7866 & tmp7879) | (tmp7866 & tmp7892) | (tmp7879 & tmp7892);
  wire tmp7894;
  assign tmp7894 = (tmp7813 & tmp7853) | (tmp7813 & tmp7893) | (tmp7853 & tmp7893);
  wire tmp7895;
  assign tmp7895 = 1'b0;
  wire tmp7896;
  assign tmp7896 = 1'b0;
  wire tmp7897;
  assign tmp7897 = 1'b0;
  wire tmp7898;
  assign tmp7898 = (tmp7895 & tmp7896) | (tmp7895 & tmp7897) | (tmp7896 & tmp7897);
  wire tmp7899;
  assign tmp7899 = 1'b0;
  wire tmp7900;
  assign tmp7900 = 1'b0;
  wire tmp7901;
  assign tmp7901 = 1'b0;
  wire tmp7902;
  assign tmp7902 = (tmp7899 & tmp7900) | (tmp7899 & tmp7901) | (tmp7900 & tmp7901);
  wire tmp7903;
  assign tmp7903 = 1'b0;
  wire tmp7904;
  assign tmp7904 = 1'b0;
  wire tmp7905;
  assign tmp7905 = 1'b0;
  wire tmp7906;
  assign tmp7906 = (tmp7903 & tmp7904) | (tmp7903 & tmp7905) | (tmp7904 & tmp7905);
  wire tmp7907;
  assign tmp7907 = (tmp7898 & tmp7902) | (tmp7898 & tmp7906) | (tmp7902 & tmp7906);
  wire tmp7908;
  assign tmp7908 = 1'b0;
  wire tmp7909;
  assign tmp7909 = 1'b0;
  wire tmp7910;
  assign tmp7910 = 1'b0;
  wire tmp7911;
  assign tmp7911 = (tmp7908 & tmp7909) | (tmp7908 & tmp7910) | (tmp7909 & tmp7910);
  wire tmp7912;
  assign tmp7912 = 1'b0;
  wire tmp7913;
  assign tmp7913 = 1'b1;
  wire tmp7914;
  assign tmp7914 = 1'b0;
  wire tmp7915;
  assign tmp7915 = (tmp7912 & tmp7913) | (tmp7912 & tmp7914) | (tmp7913 & tmp7914);
  wire tmp7916;
  assign tmp7916 = 1'b0;
  wire tmp7917;
  assign tmp7917 = 1'b0;
  wire tmp7918;
  assign tmp7918 = 1'b0;
  wire tmp7919;
  assign tmp7919 = (tmp7916 & tmp7917) | (tmp7916 & tmp7918) | (tmp7917 & tmp7918);
  wire tmp7920;
  assign tmp7920 = (tmp7911 & tmp7915) | (tmp7911 & tmp7919) | (tmp7915 & tmp7919);
  wire tmp7921;
  assign tmp7921 = 1'b0;
  wire tmp7922;
  assign tmp7922 = 1'b0;
  wire tmp7923;
  assign tmp7923 = 1'b0;
  wire tmp7924;
  assign tmp7924 = (tmp7921 & tmp7922) | (tmp7921 & tmp7923) | (tmp7922 & tmp7923);
  wire tmp7925;
  assign tmp7925 = 1'b0;
  wire tmp7926;
  assign tmp7926 = 1'b0;
  wire tmp7927;
  assign tmp7927 = 1'b0;
  wire tmp7928;
  assign tmp7928 = (tmp7925 & tmp7926) | (tmp7925 & tmp7927) | (tmp7926 & tmp7927);
  wire tmp7929;
  assign tmp7929 = 1'b0;
  wire tmp7930;
  assign tmp7930 = 1'b0;
  wire tmp7931;
  assign tmp7931 = 1'b0;
  wire tmp7932;
  assign tmp7932 = (tmp7929 & tmp7930) | (tmp7929 & tmp7931) | (tmp7930 & tmp7931);
  wire tmp7933;
  assign tmp7933 = (tmp7924 & tmp7928) | (tmp7924 & tmp7932) | (tmp7928 & tmp7932);
  wire tmp7934;
  assign tmp7934 = (tmp7907 & tmp7920) | (tmp7907 & tmp7933) | (tmp7920 & tmp7933);
  wire tmp7935;
  assign tmp7935 = 1'b0;
  wire tmp7936;
  assign tmp7936 = 1'b0;
  wire tmp7937;
  assign tmp7937 = 1'b0;
  wire tmp7938;
  assign tmp7938 = (tmp7935 & tmp7936) | (tmp7935 & tmp7937) | (tmp7936 & tmp7937);
  wire tmp7939;
  assign tmp7939 = 1'b0;
  wire tmp7940;
  assign tmp7940 = 1'b1;
  wire tmp7941;
  assign tmp7941 = 1'b0;
  wire tmp7942;
  assign tmp7942 = (tmp7939 & tmp7940) | (tmp7939 & tmp7941) | (tmp7940 & tmp7941);
  wire tmp7943;
  assign tmp7943 = 1'b0;
  wire tmp7944;
  assign tmp7944 = 1'b0;
  wire tmp7945;
  assign tmp7945 = 1'b0;
  wire tmp7946;
  assign tmp7946 = (tmp7943 & tmp7944) | (tmp7943 & tmp7945) | (tmp7944 & tmp7945);
  wire tmp7947;
  assign tmp7947 = (tmp7938 & tmp7942) | (tmp7938 & tmp7946) | (tmp7942 & tmp7946);
  wire tmp7948;
  assign tmp7948 = 1'b0;
  wire tmp7949;
  assign tmp7949 = 1'b1;
  wire tmp7950;
  assign tmp7950 = 1'b0;
  wire tmp7951;
  assign tmp7951 = (tmp7948 & tmp7949) | (tmp7948 & tmp7950) | (tmp7949 & tmp7950);
  wire tmp7952;
  assign tmp7952 = 1'b1;
  wire tmp7953;
  assign tmp7953 = ~pi6;
  wire tmp7954;
  assign tmp7954 = ~pi7;
  wire tmp7955;
  assign tmp7955 = (tmp7952 & tmp7953) | (tmp7952 & tmp7954) | (tmp7953 & tmp7954);
  wire tmp7956;
  assign tmp7956 = 1'b0;
  wire tmp7957;
  assign tmp7957 = ~pi7;
  wire tmp7958;
  assign tmp7958 = 1'b0;
  wire tmp7959;
  assign tmp7959 = (tmp7956 & tmp7957) | (tmp7956 & tmp7958) | (tmp7957 & tmp7958);
  wire tmp7960;
  assign tmp7960 = (tmp7951 & tmp7955) | (tmp7951 & tmp7959) | (tmp7955 & tmp7959);
  wire tmp7961;
  assign tmp7961 = 1'b0;
  wire tmp7962;
  assign tmp7962 = 1'b0;
  wire tmp7963;
  assign tmp7963 = 1'b0;
  wire tmp7964;
  assign tmp7964 = (tmp7961 & tmp7962) | (tmp7961 & tmp7963) | (tmp7962 & tmp7963);
  wire tmp7965;
  assign tmp7965 = 1'b0;
  wire tmp7966;
  assign tmp7966 = ~pi7;
  wire tmp7967;
  assign tmp7967 = 1'b0;
  wire tmp7968;
  assign tmp7968 = (tmp7965 & tmp7966) | (tmp7965 & tmp7967) | (tmp7966 & tmp7967);
  wire tmp7969;
  assign tmp7969 = 1'b0;
  wire tmp7970;
  assign tmp7970 = 1'b0;
  wire tmp7971;
  assign tmp7971 = 1'b0;
  wire tmp7972;
  assign tmp7972 = (tmp7969 & tmp7970) | (tmp7969 & tmp7971) | (tmp7970 & tmp7971);
  wire tmp7973;
  assign tmp7973 = (tmp7964 & tmp7968) | (tmp7964 & tmp7972) | (tmp7968 & tmp7972);
  wire tmp7974;
  assign tmp7974 = (tmp7947 & tmp7960) | (tmp7947 & tmp7973) | (tmp7960 & tmp7973);
  wire tmp7975;
  assign tmp7975 = 1'b0;
  wire tmp7976;
  assign tmp7976 = 1'b0;
  wire tmp7977;
  assign tmp7977 = 1'b0;
  wire tmp7978;
  assign tmp7978 = (tmp7975 & tmp7976) | (tmp7975 & tmp7977) | (tmp7976 & tmp7977);
  wire tmp7979;
  assign tmp7979 = 1'b0;
  wire tmp7980;
  assign tmp7980 = 1'b0;
  wire tmp7981;
  assign tmp7981 = 1'b0;
  wire tmp7982;
  assign tmp7982 = (tmp7979 & tmp7980) | (tmp7979 & tmp7981) | (tmp7980 & tmp7981);
  wire tmp7983;
  assign tmp7983 = 1'b0;
  wire tmp7984;
  assign tmp7984 = 1'b0;
  wire tmp7985;
  assign tmp7985 = 1'b0;
  wire tmp7986;
  assign tmp7986 = (tmp7983 & tmp7984) | (tmp7983 & tmp7985) | (tmp7984 & tmp7985);
  wire tmp7987;
  assign tmp7987 = (tmp7978 & tmp7982) | (tmp7978 & tmp7986) | (tmp7982 & tmp7986);
  wire tmp7988;
  assign tmp7988 = 1'b0;
  wire tmp7989;
  assign tmp7989 = 1'b0;
  wire tmp7990;
  assign tmp7990 = 1'b0;
  wire tmp7991;
  assign tmp7991 = (tmp7988 & tmp7989) | (tmp7988 & tmp7990) | (tmp7989 & tmp7990);
  wire tmp7992;
  assign tmp7992 = 1'b0;
  wire tmp7993;
  assign tmp7993 = ~pi7;
  wire tmp7994;
  assign tmp7994 = 1'b0;
  wire tmp7995;
  assign tmp7995 = (tmp7992 & tmp7993) | (tmp7992 & tmp7994) | (tmp7993 & tmp7994);
  wire tmp7996;
  assign tmp7996 = 1'b0;
  wire tmp7997;
  assign tmp7997 = 1'b0;
  wire tmp7998;
  assign tmp7998 = 1'b0;
  wire tmp7999;
  assign tmp7999 = (tmp7996 & tmp7997) | (tmp7996 & tmp7998) | (tmp7997 & tmp7998);
  wire tmp8000;
  assign tmp8000 = (tmp7991 & tmp7995) | (tmp7991 & tmp7999) | (tmp7995 & tmp7999);
  wire tmp8001;
  assign tmp8001 = 1'b0;
  wire tmp8002;
  assign tmp8002 = 1'b0;
  wire tmp8003;
  assign tmp8003 = 1'b0;
  wire tmp8004;
  assign tmp8004 = (tmp8001 & tmp8002) | (tmp8001 & tmp8003) | (tmp8002 & tmp8003);
  wire tmp8005;
  assign tmp8005 = 1'b0;
  wire tmp8006;
  assign tmp8006 = 1'b0;
  wire tmp8007;
  assign tmp8007 = 1'b0;
  wire tmp8008;
  assign tmp8008 = (tmp8005 & tmp8006) | (tmp8005 & tmp8007) | (tmp8006 & tmp8007);
  wire tmp8009;
  assign tmp8009 = 1'b0;
  wire tmp8010;
  assign tmp8010 = 1'b0;
  wire tmp8011;
  assign tmp8011 = 1'b0;
  wire tmp8012;
  assign tmp8012 = (tmp8009 & tmp8010) | (tmp8009 & tmp8011) | (tmp8010 & tmp8011);
  wire tmp8013;
  assign tmp8013 = (tmp8004 & tmp8008) | (tmp8004 & tmp8012) | (tmp8008 & tmp8012);
  wire tmp8014;
  assign tmp8014 = (tmp7987 & tmp8000) | (tmp7987 & tmp8013) | (tmp8000 & tmp8013);
  wire tmp8015;
  assign tmp8015 = (tmp7934 & tmp7974) | (tmp7934 & tmp8014) | (tmp7974 & tmp8014);
  wire tmp8016;
  assign tmp8016 = (tmp7773 & tmp7894) | (tmp7773 & tmp8015) | (tmp7894 & tmp8015);
  wire tmp8017;
  assign tmp8017 = 1'b0;
  wire tmp8018;
  assign tmp8018 = 1'b0;
  wire tmp8019;
  assign tmp8019 = 1'b0;
  wire tmp8020;
  assign tmp8020 = (tmp8017 & tmp8018) | (tmp8017 & tmp8019) | (tmp8018 & tmp8019);
  wire tmp8021;
  assign tmp8021 = 1'b0;
  wire tmp8022;
  assign tmp8022 = 1'b1;
  wire tmp8023;
  assign tmp8023 = 1'b0;
  wire tmp8024;
  assign tmp8024 = (tmp8021 & tmp8022) | (tmp8021 & tmp8023) | (tmp8022 & tmp8023);
  wire tmp8025;
  assign tmp8025 = 1'b0;
  wire tmp8026;
  assign tmp8026 = 1'b0;
  wire tmp8027;
  assign tmp8027 = 1'b0;
  wire tmp8028;
  assign tmp8028 = (tmp8025 & tmp8026) | (tmp8025 & tmp8027) | (tmp8026 & tmp8027);
  wire tmp8029;
  assign tmp8029 = (tmp8020 & tmp8024) | (tmp8020 & tmp8028) | (tmp8024 & tmp8028);
  wire tmp8030;
  assign tmp8030 = 1'b0;
  wire tmp8031;
  assign tmp8031 = 1'b1;
  wire tmp8032;
  assign tmp8032 = 1'b0;
  wire tmp8033;
  assign tmp8033 = (tmp8030 & tmp8031) | (tmp8030 & tmp8032) | (tmp8031 & tmp8032);
  wire tmp8034;
  assign tmp8034 = 1'b1;
  wire tmp8035;
  assign tmp8035 = 1'b1;
  wire tmp8036;
  assign tmp8036 = 1'b1;
  wire tmp8037;
  assign tmp8037 = (tmp8034 & tmp8035) | (tmp8034 & tmp8036) | (tmp8035 & tmp8036);
  wire tmp8038;
  assign tmp8038 = 1'b0;
  wire tmp8039;
  assign tmp8039 = 1'b1;
  wire tmp8040;
  assign tmp8040 = 1'b0;
  wire tmp8041;
  assign tmp8041 = (tmp8038 & tmp8039) | (tmp8038 & tmp8040) | (tmp8039 & tmp8040);
  wire tmp8042;
  assign tmp8042 = (tmp8033 & tmp8037) | (tmp8033 & tmp8041) | (tmp8037 & tmp8041);
  wire tmp8043;
  assign tmp8043 = 1'b0;
  wire tmp8044;
  assign tmp8044 = 1'b0;
  wire tmp8045;
  assign tmp8045 = 1'b0;
  wire tmp8046;
  assign tmp8046 = (tmp8043 & tmp8044) | (tmp8043 & tmp8045) | (tmp8044 & tmp8045);
  wire tmp8047;
  assign tmp8047 = 1'b0;
  wire tmp8048;
  assign tmp8048 = 1'b1;
  wire tmp8049;
  assign tmp8049 = 1'b0;
  wire tmp8050;
  assign tmp8050 = (tmp8047 & tmp8048) | (tmp8047 & tmp8049) | (tmp8048 & tmp8049);
  wire tmp8051;
  assign tmp8051 = 1'b0;
  wire tmp8052;
  assign tmp8052 = 1'b0;
  wire tmp8053;
  assign tmp8053 = 1'b0;
  wire tmp8054;
  assign tmp8054 = (tmp8051 & tmp8052) | (tmp8051 & tmp8053) | (tmp8052 & tmp8053);
  wire tmp8055;
  assign tmp8055 = (tmp8046 & tmp8050) | (tmp8046 & tmp8054) | (tmp8050 & tmp8054);
  wire tmp8056;
  assign tmp8056 = (tmp8029 & tmp8042) | (tmp8029 & tmp8055) | (tmp8042 & tmp8055);
  wire tmp8057;
  assign tmp8057 = 1'b0;
  wire tmp8058;
  assign tmp8058 = 1'b1;
  wire tmp8059;
  assign tmp8059 = 1'b0;
  wire tmp8060;
  assign tmp8060 = (tmp8057 & tmp8058) | (tmp8057 & tmp8059) | (tmp8058 & tmp8059);
  wire tmp8061;
  assign tmp8061 = 1'b1;
  wire tmp8062;
  assign tmp8062 = 1'b1;
  wire tmp8063;
  assign tmp8063 = 1'b1;
  wire tmp8064;
  assign tmp8064 = (tmp8061 & tmp8062) | (tmp8061 & tmp8063) | (tmp8062 & tmp8063);
  wire tmp8065;
  assign tmp8065 = 1'b0;
  wire tmp8066;
  assign tmp8066 = 1'b1;
  wire tmp8067;
  assign tmp8067 = 1'b0;
  wire tmp8068;
  assign tmp8068 = (tmp8065 & tmp8066) | (tmp8065 & tmp8067) | (tmp8066 & tmp8067);
  wire tmp8069;
  assign tmp8069 = (tmp8060 & tmp8064) | (tmp8060 & tmp8068) | (tmp8064 & tmp8068);
  wire tmp8070;
  assign tmp8070 = 1'b1;
  wire tmp8071;
  assign tmp8071 = 1'b1;
  wire tmp8072;
  assign tmp8072 = 1'b1;
  wire tmp8073;
  assign tmp8073 = (tmp8070 & tmp8071) | (tmp8070 & tmp8072) | (tmp8071 & tmp8072);
  wire tmp8074;
  assign tmp8074 = 1'b1;
  wire tmp8075;
  assign tmp8075 = ~pi5;
  wire tmp8076;
  assign tmp8076 = ~pi6;
  wire tmp8077;
  assign tmp8077 = (tmp8074 & tmp8075) | (tmp8074 & tmp8076) | (tmp8075 & tmp8076);
  wire tmp8078;
  assign tmp8078 = 1'b1;
  wire tmp8079;
  assign tmp8079 = ~pi6;
  wire tmp8080;
  assign tmp8080 = ~pi7;
  wire tmp8081;
  assign tmp8081 = (tmp8078 & tmp8079) | (tmp8078 & tmp8080) | (tmp8079 & tmp8080);
  wire tmp8082;
  assign tmp8082 = (tmp8073 & tmp8077) | (tmp8073 & tmp8081) | (tmp8077 & tmp8081);
  wire tmp8083;
  assign tmp8083 = 1'b0;
  wire tmp8084;
  assign tmp8084 = 1'b1;
  wire tmp8085;
  assign tmp8085 = 1'b0;
  wire tmp8086;
  assign tmp8086 = (tmp8083 & tmp8084) | (tmp8083 & tmp8085) | (tmp8084 & tmp8085);
  wire tmp8087;
  assign tmp8087 = 1'b1;
  wire tmp8088;
  assign tmp8088 = ~pi6;
  wire tmp8089;
  assign tmp8089 = ~pi7;
  wire tmp8090;
  assign tmp8090 = (tmp8087 & tmp8088) | (tmp8087 & tmp8089) | (tmp8088 & tmp8089);
  wire tmp8091;
  assign tmp8091 = 1'b0;
  wire tmp8092;
  assign tmp8092 = ~pi7;
  wire tmp8093;
  assign tmp8093 = 1'b0;
  wire tmp8094;
  assign tmp8094 = (tmp8091 & tmp8092) | (tmp8091 & tmp8093) | (tmp8092 & tmp8093);
  wire tmp8095;
  assign tmp8095 = (tmp8086 & tmp8090) | (tmp8086 & tmp8094) | (tmp8090 & tmp8094);
  wire tmp8096;
  assign tmp8096 = (tmp8069 & tmp8082) | (tmp8069 & tmp8095) | (tmp8082 & tmp8095);
  wire tmp8097;
  assign tmp8097 = 1'b0;
  wire tmp8098;
  assign tmp8098 = 1'b0;
  wire tmp8099;
  assign tmp8099 = 1'b0;
  wire tmp8100;
  assign tmp8100 = (tmp8097 & tmp8098) | (tmp8097 & tmp8099) | (tmp8098 & tmp8099);
  wire tmp8101;
  assign tmp8101 = 1'b0;
  wire tmp8102;
  assign tmp8102 = 1'b1;
  wire tmp8103;
  assign tmp8103 = 1'b0;
  wire tmp8104;
  assign tmp8104 = (tmp8101 & tmp8102) | (tmp8101 & tmp8103) | (tmp8102 & tmp8103);
  wire tmp8105;
  assign tmp8105 = 1'b0;
  wire tmp8106;
  assign tmp8106 = 1'b0;
  wire tmp8107;
  assign tmp8107 = 1'b0;
  wire tmp8108;
  assign tmp8108 = (tmp8105 & tmp8106) | (tmp8105 & tmp8107) | (tmp8106 & tmp8107);
  wire tmp8109;
  assign tmp8109 = (tmp8100 & tmp8104) | (tmp8100 & tmp8108) | (tmp8104 & tmp8108);
  wire tmp8110;
  assign tmp8110 = 1'b0;
  wire tmp8111;
  assign tmp8111 = 1'b1;
  wire tmp8112;
  assign tmp8112 = 1'b0;
  wire tmp8113;
  assign tmp8113 = (tmp8110 & tmp8111) | (tmp8110 & tmp8112) | (tmp8111 & tmp8112);
  wire tmp8114;
  assign tmp8114 = 1'b1;
  wire tmp8115;
  assign tmp8115 = ~pi6;
  wire tmp8116;
  assign tmp8116 = ~pi7;
  wire tmp8117;
  assign tmp8117 = (tmp8114 & tmp8115) | (tmp8114 & tmp8116) | (tmp8115 & tmp8116);
  wire tmp8118;
  assign tmp8118 = 1'b0;
  wire tmp8119;
  assign tmp8119 = ~pi7;
  wire tmp8120;
  assign tmp8120 = 1'b0;
  wire tmp8121;
  assign tmp8121 = (tmp8118 & tmp8119) | (tmp8118 & tmp8120) | (tmp8119 & tmp8120);
  wire tmp8122;
  assign tmp8122 = (tmp8113 & tmp8117) | (tmp8113 & tmp8121) | (tmp8117 & tmp8121);
  wire tmp8123;
  assign tmp8123 = 1'b0;
  wire tmp8124;
  assign tmp8124 = 1'b0;
  wire tmp8125;
  assign tmp8125 = 1'b0;
  wire tmp8126;
  assign tmp8126 = (tmp8123 & tmp8124) | (tmp8123 & tmp8125) | (tmp8124 & tmp8125);
  wire tmp8127;
  assign tmp8127 = 1'b0;
  wire tmp8128;
  assign tmp8128 = ~pi7;
  wire tmp8129;
  assign tmp8129 = 1'b0;
  wire tmp8130;
  assign tmp8130 = (tmp8127 & tmp8128) | (tmp8127 & tmp8129) | (tmp8128 & tmp8129);
  wire tmp8131;
  assign tmp8131 = 1'b0;
  wire tmp8132;
  assign tmp8132 = 1'b0;
  wire tmp8133;
  assign tmp8133 = 1'b0;
  wire tmp8134;
  assign tmp8134 = (tmp8131 & tmp8132) | (tmp8131 & tmp8133) | (tmp8132 & tmp8133);
  wire tmp8135;
  assign tmp8135 = (tmp8126 & tmp8130) | (tmp8126 & tmp8134) | (tmp8130 & tmp8134);
  wire tmp8136;
  assign tmp8136 = (tmp8109 & tmp8122) | (tmp8109 & tmp8135) | (tmp8122 & tmp8135);
  wire tmp8137;
  assign tmp8137 = (tmp8056 & tmp8096) | (tmp8056 & tmp8136) | (tmp8096 & tmp8136);
  wire tmp8138;
  assign tmp8138 = 1'b0;
  wire tmp8139;
  assign tmp8139 = 1'b1;
  wire tmp8140;
  assign tmp8140 = 1'b0;
  wire tmp8141;
  assign tmp8141 = (tmp8138 & tmp8139) | (tmp8138 & tmp8140) | (tmp8139 & tmp8140);
  wire tmp8142;
  assign tmp8142 = 1'b1;
  wire tmp8143;
  assign tmp8143 = 1'b1;
  wire tmp8144;
  assign tmp8144 = 1'b1;
  wire tmp8145;
  assign tmp8145 = (tmp8142 & tmp8143) | (tmp8142 & tmp8144) | (tmp8143 & tmp8144);
  wire tmp8146;
  assign tmp8146 = 1'b0;
  wire tmp8147;
  assign tmp8147 = 1'b1;
  wire tmp8148;
  assign tmp8148 = 1'b0;
  wire tmp8149;
  assign tmp8149 = (tmp8146 & tmp8147) | (tmp8146 & tmp8148) | (tmp8147 & tmp8148);
  wire tmp8150;
  assign tmp8150 = (tmp8141 & tmp8145) | (tmp8141 & tmp8149) | (tmp8145 & tmp8149);
  wire tmp8151;
  assign tmp8151 = 1'b1;
  wire tmp8152;
  assign tmp8152 = 1'b1;
  wire tmp8153;
  assign tmp8153 = 1'b1;
  wire tmp8154;
  assign tmp8154 = (tmp8151 & tmp8152) | (tmp8151 & tmp8153) | (tmp8152 & tmp8153);
  wire tmp8155;
  assign tmp8155 = 1'b1;
  wire tmp8156;
  assign tmp8156 = ~pi5;
  wire tmp8157;
  assign tmp8157 = ~pi6;
  wire tmp8158;
  assign tmp8158 = (tmp8155 & tmp8156) | (tmp8155 & tmp8157) | (tmp8156 & tmp8157);
  wire tmp8159;
  assign tmp8159 = 1'b1;
  wire tmp8160;
  assign tmp8160 = ~pi6;
  wire tmp8161;
  assign tmp8161 = ~pi7;
  wire tmp8162;
  assign tmp8162 = (tmp8159 & tmp8160) | (tmp8159 & tmp8161) | (tmp8160 & tmp8161);
  wire tmp8163;
  assign tmp8163 = (tmp8154 & tmp8158) | (tmp8154 & tmp8162) | (tmp8158 & tmp8162);
  wire tmp8164;
  assign tmp8164 = 1'b0;
  wire tmp8165;
  assign tmp8165 = 1'b1;
  wire tmp8166;
  assign tmp8166 = 1'b0;
  wire tmp8167;
  assign tmp8167 = (tmp8164 & tmp8165) | (tmp8164 & tmp8166) | (tmp8165 & tmp8166);
  wire tmp8168;
  assign tmp8168 = 1'b1;
  wire tmp8169;
  assign tmp8169 = ~pi6;
  wire tmp8170;
  assign tmp8170 = ~pi7;
  wire tmp8171;
  assign tmp8171 = (tmp8168 & tmp8169) | (tmp8168 & tmp8170) | (tmp8169 & tmp8170);
  wire tmp8172;
  assign tmp8172 = 1'b0;
  wire tmp8173;
  assign tmp8173 = ~pi7;
  wire tmp8174;
  assign tmp8174 = 1'b0;
  wire tmp8175;
  assign tmp8175 = (tmp8172 & tmp8173) | (tmp8172 & tmp8174) | (tmp8173 & tmp8174);
  wire tmp8176;
  assign tmp8176 = (tmp8167 & tmp8171) | (tmp8167 & tmp8175) | (tmp8171 & tmp8175);
  wire tmp8177;
  assign tmp8177 = (tmp8150 & tmp8163) | (tmp8150 & tmp8176) | (tmp8163 & tmp8176);
  wire tmp8178;
  assign tmp8178 = 1'b1;
  wire tmp8179;
  assign tmp8179 = 1'b1;
  wire tmp8180;
  assign tmp8180 = 1'b1;
  wire tmp8181;
  assign tmp8181 = (tmp8178 & tmp8179) | (tmp8178 & tmp8180) | (tmp8179 & tmp8180);
  wire tmp8182;
  assign tmp8182 = 1'b1;
  wire tmp8183;
  assign tmp8183 = ~pi5;
  wire tmp8184;
  assign tmp8184 = ~pi6;
  wire tmp8185;
  assign tmp8185 = (tmp8182 & tmp8183) | (tmp8182 & tmp8184) | (tmp8183 & tmp8184);
  wire tmp8186;
  assign tmp8186 = 1'b1;
  wire tmp8187;
  assign tmp8187 = ~pi6;
  wire tmp8188;
  assign tmp8188 = ~pi7;
  wire tmp8189;
  assign tmp8189 = (tmp8186 & tmp8187) | (tmp8186 & tmp8188) | (tmp8187 & tmp8188);
  wire tmp8190;
  assign tmp8190 = (tmp8181 & tmp8185) | (tmp8181 & tmp8189) | (tmp8185 & tmp8189);
  wire tmp8191;
  assign tmp8191 = 1'b1;
  wire tmp8192;
  assign tmp8192 = ~pi5;
  wire tmp8193;
  assign tmp8193 = ~pi6;
  wire tmp8194;
  assign tmp8194 = (tmp8191 & tmp8192) | (tmp8191 & tmp8193) | (tmp8192 & tmp8193);
  wire tmp8195;
  assign tmp8195 = ~pi5;
  wire tmp8196;
  assign tmp8196 = 1'b1;
  wire tmp8197;
  assign tmp8197 = 1'b1;
  wire tmp8198;
  assign tmp8198 = (tmp8195 & tmp8196) | (tmp8195 & tmp8197) | (tmp8196 & tmp8197);
  wire tmp8199;
  assign tmp8199 = ~pi6;
  wire tmp8200;
  assign tmp8200 = 1'b1;
  wire tmp8201;
  assign tmp8201 = 1'b1;
  wire tmp8202;
  assign tmp8202 = (tmp8199 & tmp8200) | (tmp8199 & tmp8201) | (tmp8200 & tmp8201);
  wire tmp8203;
  assign tmp8203 = (tmp8194 & tmp8198) | (tmp8194 & tmp8202) | (tmp8198 & tmp8202);
  wire tmp8204;
  assign tmp8204 = 1'b1;
  wire tmp8205;
  assign tmp8205 = ~pi6;
  wire tmp8206;
  assign tmp8206 = ~pi7;
  wire tmp8207;
  assign tmp8207 = (tmp8204 & tmp8205) | (tmp8204 & tmp8206) | (tmp8205 & tmp8206);
  wire tmp8208;
  assign tmp8208 = ~pi6;
  wire tmp8209;
  assign tmp8209 = 1'b1;
  wire tmp8210;
  assign tmp8210 = 1'b1;
  wire tmp8211;
  assign tmp8211 = (tmp8208 & tmp8209) | (tmp8208 & tmp8210) | (tmp8209 & tmp8210);
  wire tmp8212;
  assign tmp8212 = ~pi7;
  wire tmp8213;
  assign tmp8213 = 1'b1;
  wire tmp8214;
  assign tmp8214 = 1'b0;
  wire tmp8215;
  assign tmp8215 = (tmp8212 & tmp8213) | (tmp8212 & tmp8214) | (tmp8213 & tmp8214);
  wire tmp8216;
  assign tmp8216 = (tmp8207 & tmp8211) | (tmp8207 & tmp8215) | (tmp8211 & tmp8215);
  wire tmp8217;
  assign tmp8217 = (tmp8190 & tmp8203) | (tmp8190 & tmp8216) | (tmp8203 & tmp8216);
  wire tmp8218;
  assign tmp8218 = 1'b0;
  wire tmp8219;
  assign tmp8219 = 1'b1;
  wire tmp8220;
  assign tmp8220 = 1'b0;
  wire tmp8221;
  assign tmp8221 = (tmp8218 & tmp8219) | (tmp8218 & tmp8220) | (tmp8219 & tmp8220);
  wire tmp8222;
  assign tmp8222 = 1'b1;
  wire tmp8223;
  assign tmp8223 = ~pi6;
  wire tmp8224;
  assign tmp8224 = ~pi7;
  wire tmp8225;
  assign tmp8225 = (tmp8222 & tmp8223) | (tmp8222 & tmp8224) | (tmp8223 & tmp8224);
  wire tmp8226;
  assign tmp8226 = 1'b0;
  wire tmp8227;
  assign tmp8227 = ~pi7;
  wire tmp8228;
  assign tmp8228 = 1'b0;
  wire tmp8229;
  assign tmp8229 = (tmp8226 & tmp8227) | (tmp8226 & tmp8228) | (tmp8227 & tmp8228);
  wire tmp8230;
  assign tmp8230 = (tmp8221 & tmp8225) | (tmp8221 & tmp8229) | (tmp8225 & tmp8229);
  wire tmp8231;
  assign tmp8231 = 1'b1;
  wire tmp8232;
  assign tmp8232 = ~pi6;
  wire tmp8233;
  assign tmp8233 = ~pi7;
  wire tmp8234;
  assign tmp8234 = (tmp8231 & tmp8232) | (tmp8231 & tmp8233) | (tmp8232 & tmp8233);
  wire tmp8235;
  assign tmp8235 = ~pi6;
  wire tmp8236;
  assign tmp8236 = 1'b1;
  wire tmp8237;
  assign tmp8237 = 1'b1;
  wire tmp8238;
  assign tmp8238 = (tmp8235 & tmp8236) | (tmp8235 & tmp8237) | (tmp8236 & tmp8237);
  wire tmp8239;
  assign tmp8239 = ~pi7;
  wire tmp8240;
  assign tmp8240 = 1'b1;
  wire tmp8241;
  assign tmp8241 = 1'b0;
  wire tmp8242;
  assign tmp8242 = (tmp8239 & tmp8240) | (tmp8239 & tmp8241) | (tmp8240 & tmp8241);
  wire tmp8243;
  assign tmp8243 = (tmp8234 & tmp8238) | (tmp8234 & tmp8242) | (tmp8238 & tmp8242);
  wire tmp8244;
  assign tmp8244 = 1'b0;
  wire tmp8245;
  assign tmp8245 = ~pi7;
  wire tmp8246;
  assign tmp8246 = 1'b0;
  wire tmp8247;
  assign tmp8247 = (tmp8244 & tmp8245) | (tmp8244 & tmp8246) | (tmp8245 & tmp8246);
  wire tmp8248;
  assign tmp8248 = ~pi7;
  wire tmp8249;
  assign tmp8249 = 1'b1;
  wire tmp8250;
  assign tmp8250 = 1'b0;
  wire tmp8251;
  assign tmp8251 = (tmp8248 & tmp8249) | (tmp8248 & tmp8250) | (tmp8249 & tmp8250);
  wire tmp8252;
  assign tmp8252 = 1'b0;
  wire tmp8253;
  assign tmp8253 = 1'b0;
  wire tmp8254;
  assign tmp8254 = 1'b0;
  wire tmp8255;
  assign tmp8255 = (tmp8252 & tmp8253) | (tmp8252 & tmp8254) | (tmp8253 & tmp8254);
  wire tmp8256;
  assign tmp8256 = (tmp8247 & tmp8251) | (tmp8247 & tmp8255) | (tmp8251 & tmp8255);
  wire tmp8257;
  assign tmp8257 = (tmp8230 & tmp8243) | (tmp8230 & tmp8256) | (tmp8243 & tmp8256);
  wire tmp8258;
  assign tmp8258 = (tmp8177 & tmp8217) | (tmp8177 & tmp8257) | (tmp8217 & tmp8257);
  wire tmp8259;
  assign tmp8259 = 1'b0;
  wire tmp8260;
  assign tmp8260 = 1'b0;
  wire tmp8261;
  assign tmp8261 = 1'b0;
  wire tmp8262;
  assign tmp8262 = (tmp8259 & tmp8260) | (tmp8259 & tmp8261) | (tmp8260 & tmp8261);
  wire tmp8263;
  assign tmp8263 = 1'b0;
  wire tmp8264;
  assign tmp8264 = 1'b1;
  wire tmp8265;
  assign tmp8265 = 1'b0;
  wire tmp8266;
  assign tmp8266 = (tmp8263 & tmp8264) | (tmp8263 & tmp8265) | (tmp8264 & tmp8265);
  wire tmp8267;
  assign tmp8267 = 1'b0;
  wire tmp8268;
  assign tmp8268 = 1'b0;
  wire tmp8269;
  assign tmp8269 = 1'b0;
  wire tmp8270;
  assign tmp8270 = (tmp8267 & tmp8268) | (tmp8267 & tmp8269) | (tmp8268 & tmp8269);
  wire tmp8271;
  assign tmp8271 = (tmp8262 & tmp8266) | (tmp8262 & tmp8270) | (tmp8266 & tmp8270);
  wire tmp8272;
  assign tmp8272 = 1'b0;
  wire tmp8273;
  assign tmp8273 = 1'b1;
  wire tmp8274;
  assign tmp8274 = 1'b0;
  wire tmp8275;
  assign tmp8275 = (tmp8272 & tmp8273) | (tmp8272 & tmp8274) | (tmp8273 & tmp8274);
  wire tmp8276;
  assign tmp8276 = 1'b1;
  wire tmp8277;
  assign tmp8277 = ~pi6;
  wire tmp8278;
  assign tmp8278 = ~pi7;
  wire tmp8279;
  assign tmp8279 = (tmp8276 & tmp8277) | (tmp8276 & tmp8278) | (tmp8277 & tmp8278);
  wire tmp8280;
  assign tmp8280 = 1'b0;
  wire tmp8281;
  assign tmp8281 = ~pi7;
  wire tmp8282;
  assign tmp8282 = 1'b0;
  wire tmp8283;
  assign tmp8283 = (tmp8280 & tmp8281) | (tmp8280 & tmp8282) | (tmp8281 & tmp8282);
  wire tmp8284;
  assign tmp8284 = (tmp8275 & tmp8279) | (tmp8275 & tmp8283) | (tmp8279 & tmp8283);
  wire tmp8285;
  assign tmp8285 = 1'b0;
  wire tmp8286;
  assign tmp8286 = 1'b0;
  wire tmp8287;
  assign tmp8287 = 1'b0;
  wire tmp8288;
  assign tmp8288 = (tmp8285 & tmp8286) | (tmp8285 & tmp8287) | (tmp8286 & tmp8287);
  wire tmp8289;
  assign tmp8289 = 1'b0;
  wire tmp8290;
  assign tmp8290 = ~pi7;
  wire tmp8291;
  assign tmp8291 = 1'b0;
  wire tmp8292;
  assign tmp8292 = (tmp8289 & tmp8290) | (tmp8289 & tmp8291) | (tmp8290 & tmp8291);
  wire tmp8293;
  assign tmp8293 = 1'b0;
  wire tmp8294;
  assign tmp8294 = 1'b0;
  wire tmp8295;
  assign tmp8295 = 1'b0;
  wire tmp8296;
  assign tmp8296 = (tmp8293 & tmp8294) | (tmp8293 & tmp8295) | (tmp8294 & tmp8295);
  wire tmp8297;
  assign tmp8297 = (tmp8288 & tmp8292) | (tmp8288 & tmp8296) | (tmp8292 & tmp8296);
  wire tmp8298;
  assign tmp8298 = (tmp8271 & tmp8284) | (tmp8271 & tmp8297) | (tmp8284 & tmp8297);
  wire tmp8299;
  assign tmp8299 = 1'b0;
  wire tmp8300;
  assign tmp8300 = 1'b1;
  wire tmp8301;
  assign tmp8301 = 1'b0;
  wire tmp8302;
  assign tmp8302 = (tmp8299 & tmp8300) | (tmp8299 & tmp8301) | (tmp8300 & tmp8301);
  wire tmp8303;
  assign tmp8303 = 1'b1;
  wire tmp8304;
  assign tmp8304 = ~pi6;
  wire tmp8305;
  assign tmp8305 = ~pi7;
  wire tmp8306;
  assign tmp8306 = (tmp8303 & tmp8304) | (tmp8303 & tmp8305) | (tmp8304 & tmp8305);
  wire tmp8307;
  assign tmp8307 = 1'b0;
  wire tmp8308;
  assign tmp8308 = ~pi7;
  wire tmp8309;
  assign tmp8309 = 1'b0;
  wire tmp8310;
  assign tmp8310 = (tmp8307 & tmp8308) | (tmp8307 & tmp8309) | (tmp8308 & tmp8309);
  wire tmp8311;
  assign tmp8311 = (tmp8302 & tmp8306) | (tmp8302 & tmp8310) | (tmp8306 & tmp8310);
  wire tmp8312;
  assign tmp8312 = 1'b1;
  wire tmp8313;
  assign tmp8313 = ~pi6;
  wire tmp8314;
  assign tmp8314 = ~pi7;
  wire tmp8315;
  assign tmp8315 = (tmp8312 & tmp8313) | (tmp8312 & tmp8314) | (tmp8313 & tmp8314);
  wire tmp8316;
  assign tmp8316 = ~pi6;
  wire tmp8317;
  assign tmp8317 = 1'b1;
  wire tmp8318;
  assign tmp8318 = 1'b1;
  wire tmp8319;
  assign tmp8319 = (tmp8316 & tmp8317) | (tmp8316 & tmp8318) | (tmp8317 & tmp8318);
  wire tmp8320;
  assign tmp8320 = ~pi7;
  wire tmp8321;
  assign tmp8321 = 1'b1;
  wire tmp8322;
  assign tmp8322 = 1'b0;
  wire tmp8323;
  assign tmp8323 = (tmp8320 & tmp8321) | (tmp8320 & tmp8322) | (tmp8321 & tmp8322);
  wire tmp8324;
  assign tmp8324 = (tmp8315 & tmp8319) | (tmp8315 & tmp8323) | (tmp8319 & tmp8323);
  wire tmp8325;
  assign tmp8325 = 1'b0;
  wire tmp8326;
  assign tmp8326 = ~pi7;
  wire tmp8327;
  assign tmp8327 = 1'b0;
  wire tmp8328;
  assign tmp8328 = (tmp8325 & tmp8326) | (tmp8325 & tmp8327) | (tmp8326 & tmp8327);
  wire tmp8329;
  assign tmp8329 = ~pi7;
  wire tmp8330;
  assign tmp8330 = 1'b1;
  wire tmp8331;
  assign tmp8331 = 1'b0;
  wire tmp8332;
  assign tmp8332 = (tmp8329 & tmp8330) | (tmp8329 & tmp8331) | (tmp8330 & tmp8331);
  wire tmp8333;
  assign tmp8333 = 1'b0;
  wire tmp8334;
  assign tmp8334 = 1'b0;
  wire tmp8335;
  assign tmp8335 = 1'b0;
  wire tmp8336;
  assign tmp8336 = (tmp8333 & tmp8334) | (tmp8333 & tmp8335) | (tmp8334 & tmp8335);
  wire tmp8337;
  assign tmp8337 = (tmp8328 & tmp8332) | (tmp8328 & tmp8336) | (tmp8332 & tmp8336);
  wire tmp8338;
  assign tmp8338 = (tmp8311 & tmp8324) | (tmp8311 & tmp8337) | (tmp8324 & tmp8337);
  wire tmp8339;
  assign tmp8339 = 1'b0;
  wire tmp8340;
  assign tmp8340 = 1'b0;
  wire tmp8341;
  assign tmp8341 = 1'b0;
  wire tmp8342;
  assign tmp8342 = (tmp8339 & tmp8340) | (tmp8339 & tmp8341) | (tmp8340 & tmp8341);
  wire tmp8343;
  assign tmp8343 = 1'b0;
  wire tmp8344;
  assign tmp8344 = ~pi7;
  wire tmp8345;
  assign tmp8345 = 1'b0;
  wire tmp8346;
  assign tmp8346 = (tmp8343 & tmp8344) | (tmp8343 & tmp8345) | (tmp8344 & tmp8345);
  wire tmp8347;
  assign tmp8347 = 1'b0;
  wire tmp8348;
  assign tmp8348 = 1'b0;
  wire tmp8349;
  assign tmp8349 = 1'b0;
  wire tmp8350;
  assign tmp8350 = (tmp8347 & tmp8348) | (tmp8347 & tmp8349) | (tmp8348 & tmp8349);
  wire tmp8351;
  assign tmp8351 = (tmp8342 & tmp8346) | (tmp8342 & tmp8350) | (tmp8346 & tmp8350);
  wire tmp8352;
  assign tmp8352 = 1'b0;
  wire tmp8353;
  assign tmp8353 = ~pi7;
  wire tmp8354;
  assign tmp8354 = 1'b0;
  wire tmp8355;
  assign tmp8355 = (tmp8352 & tmp8353) | (tmp8352 & tmp8354) | (tmp8353 & tmp8354);
  wire tmp8356;
  assign tmp8356 = ~pi7;
  wire tmp8357;
  assign tmp8357 = 1'b1;
  wire tmp8358;
  assign tmp8358 = 1'b0;
  wire tmp8359;
  assign tmp8359 = (tmp8356 & tmp8357) | (tmp8356 & tmp8358) | (tmp8357 & tmp8358);
  wire tmp8360;
  assign tmp8360 = 1'b0;
  wire tmp8361;
  assign tmp8361 = 1'b0;
  wire tmp8362;
  assign tmp8362 = 1'b0;
  wire tmp8363;
  assign tmp8363 = (tmp8360 & tmp8361) | (tmp8360 & tmp8362) | (tmp8361 & tmp8362);
  wire tmp8364;
  assign tmp8364 = (tmp8355 & tmp8359) | (tmp8355 & tmp8363) | (tmp8359 & tmp8363);
  wire tmp8365;
  assign tmp8365 = 1'b0;
  wire tmp8366;
  assign tmp8366 = 1'b0;
  wire tmp8367;
  assign tmp8367 = 1'b0;
  wire tmp8368;
  assign tmp8368 = (tmp8365 & tmp8366) | (tmp8365 & tmp8367) | (tmp8366 & tmp8367);
  wire tmp8369;
  assign tmp8369 = 1'b0;
  wire tmp8370;
  assign tmp8370 = 1'b0;
  wire tmp8371;
  assign tmp8371 = 1'b0;
  wire tmp8372;
  assign tmp8372 = (tmp8369 & tmp8370) | (tmp8369 & tmp8371) | (tmp8370 & tmp8371);
  wire tmp8373;
  assign tmp8373 = 1'b0;
  wire tmp8374;
  assign tmp8374 = 1'b0;
  wire tmp8375;
  assign tmp8375 = 1'b0;
  wire tmp8376;
  assign tmp8376 = (tmp8373 & tmp8374) | (tmp8373 & tmp8375) | (tmp8374 & tmp8375);
  wire tmp8377;
  assign tmp8377 = (tmp8368 & tmp8372) | (tmp8368 & tmp8376) | (tmp8372 & tmp8376);
  wire tmp8378;
  assign tmp8378 = (tmp8351 & tmp8364) | (tmp8351 & tmp8377) | (tmp8364 & tmp8377);
  wire tmp8379;
  assign tmp8379 = (tmp8298 & tmp8338) | (tmp8298 & tmp8378) | (tmp8338 & tmp8378);
  wire tmp8380;
  assign tmp8380 = (tmp8137 & tmp8258) | (tmp8137 & tmp8379) | (tmp8258 & tmp8379);
  wire tmp8381;
  assign tmp8381 = 1'b0;
  wire tmp8382;
  assign tmp8382 = 1'b0;
  wire tmp8383;
  assign tmp8383 = 1'b0;
  wire tmp8384;
  assign tmp8384 = (tmp8381 & tmp8382) | (tmp8381 & tmp8383) | (tmp8382 & tmp8383);
  wire tmp8385;
  assign tmp8385 = 1'b0;
  wire tmp8386;
  assign tmp8386 = 1'b0;
  wire tmp8387;
  assign tmp8387 = 1'b0;
  wire tmp8388;
  assign tmp8388 = (tmp8385 & tmp8386) | (tmp8385 & tmp8387) | (tmp8386 & tmp8387);
  wire tmp8389;
  assign tmp8389 = 1'b0;
  wire tmp8390;
  assign tmp8390 = 1'b0;
  wire tmp8391;
  assign tmp8391 = 1'b0;
  wire tmp8392;
  assign tmp8392 = (tmp8389 & tmp8390) | (tmp8389 & tmp8391) | (tmp8390 & tmp8391);
  wire tmp8393;
  assign tmp8393 = (tmp8384 & tmp8388) | (tmp8384 & tmp8392) | (tmp8388 & tmp8392);
  wire tmp8394;
  assign tmp8394 = 1'b0;
  wire tmp8395;
  assign tmp8395 = 1'b0;
  wire tmp8396;
  assign tmp8396 = 1'b0;
  wire tmp8397;
  assign tmp8397 = (tmp8394 & tmp8395) | (tmp8394 & tmp8396) | (tmp8395 & tmp8396);
  wire tmp8398;
  assign tmp8398 = 1'b0;
  wire tmp8399;
  assign tmp8399 = 1'b1;
  wire tmp8400;
  assign tmp8400 = 1'b0;
  wire tmp8401;
  assign tmp8401 = (tmp8398 & tmp8399) | (tmp8398 & tmp8400) | (tmp8399 & tmp8400);
  wire tmp8402;
  assign tmp8402 = 1'b0;
  wire tmp8403;
  assign tmp8403 = 1'b0;
  wire tmp8404;
  assign tmp8404 = 1'b0;
  wire tmp8405;
  assign tmp8405 = (tmp8402 & tmp8403) | (tmp8402 & tmp8404) | (tmp8403 & tmp8404);
  wire tmp8406;
  assign tmp8406 = (tmp8397 & tmp8401) | (tmp8397 & tmp8405) | (tmp8401 & tmp8405);
  wire tmp8407;
  assign tmp8407 = 1'b0;
  wire tmp8408;
  assign tmp8408 = 1'b0;
  wire tmp8409;
  assign tmp8409 = 1'b0;
  wire tmp8410;
  assign tmp8410 = (tmp8407 & tmp8408) | (tmp8407 & tmp8409) | (tmp8408 & tmp8409);
  wire tmp8411;
  assign tmp8411 = 1'b0;
  wire tmp8412;
  assign tmp8412 = 1'b0;
  wire tmp8413;
  assign tmp8413 = 1'b0;
  wire tmp8414;
  assign tmp8414 = (tmp8411 & tmp8412) | (tmp8411 & tmp8413) | (tmp8412 & tmp8413);
  wire tmp8415;
  assign tmp8415 = 1'b0;
  wire tmp8416;
  assign tmp8416 = 1'b0;
  wire tmp8417;
  assign tmp8417 = 1'b0;
  wire tmp8418;
  assign tmp8418 = (tmp8415 & tmp8416) | (tmp8415 & tmp8417) | (tmp8416 & tmp8417);
  wire tmp8419;
  assign tmp8419 = (tmp8410 & tmp8414) | (tmp8410 & tmp8418) | (tmp8414 & tmp8418);
  wire tmp8420;
  assign tmp8420 = (tmp8393 & tmp8406) | (tmp8393 & tmp8419) | (tmp8406 & tmp8419);
  wire tmp8421;
  assign tmp8421 = 1'b0;
  wire tmp8422;
  assign tmp8422 = 1'b0;
  wire tmp8423;
  assign tmp8423 = 1'b0;
  wire tmp8424;
  assign tmp8424 = (tmp8421 & tmp8422) | (tmp8421 & tmp8423) | (tmp8422 & tmp8423);
  wire tmp8425;
  assign tmp8425 = 1'b0;
  wire tmp8426;
  assign tmp8426 = 1'b1;
  wire tmp8427;
  assign tmp8427 = 1'b0;
  wire tmp8428;
  assign tmp8428 = (tmp8425 & tmp8426) | (tmp8425 & tmp8427) | (tmp8426 & tmp8427);
  wire tmp8429;
  assign tmp8429 = 1'b0;
  wire tmp8430;
  assign tmp8430 = 1'b0;
  wire tmp8431;
  assign tmp8431 = 1'b0;
  wire tmp8432;
  assign tmp8432 = (tmp8429 & tmp8430) | (tmp8429 & tmp8431) | (tmp8430 & tmp8431);
  wire tmp8433;
  assign tmp8433 = (tmp8424 & tmp8428) | (tmp8424 & tmp8432) | (tmp8428 & tmp8432);
  wire tmp8434;
  assign tmp8434 = 1'b0;
  wire tmp8435;
  assign tmp8435 = 1'b1;
  wire tmp8436;
  assign tmp8436 = 1'b0;
  wire tmp8437;
  assign tmp8437 = (tmp8434 & tmp8435) | (tmp8434 & tmp8436) | (tmp8435 & tmp8436);
  wire tmp8438;
  assign tmp8438 = 1'b1;
  wire tmp8439;
  assign tmp8439 = ~pi6;
  wire tmp8440;
  assign tmp8440 = ~pi7;
  wire tmp8441;
  assign tmp8441 = (tmp8438 & tmp8439) | (tmp8438 & tmp8440) | (tmp8439 & tmp8440);
  wire tmp8442;
  assign tmp8442 = 1'b0;
  wire tmp8443;
  assign tmp8443 = ~pi7;
  wire tmp8444;
  assign tmp8444 = 1'b0;
  wire tmp8445;
  assign tmp8445 = (tmp8442 & tmp8443) | (tmp8442 & tmp8444) | (tmp8443 & tmp8444);
  wire tmp8446;
  assign tmp8446 = (tmp8437 & tmp8441) | (tmp8437 & tmp8445) | (tmp8441 & tmp8445);
  wire tmp8447;
  assign tmp8447 = 1'b0;
  wire tmp8448;
  assign tmp8448 = 1'b0;
  wire tmp8449;
  assign tmp8449 = 1'b0;
  wire tmp8450;
  assign tmp8450 = (tmp8447 & tmp8448) | (tmp8447 & tmp8449) | (tmp8448 & tmp8449);
  wire tmp8451;
  assign tmp8451 = 1'b0;
  wire tmp8452;
  assign tmp8452 = ~pi7;
  wire tmp8453;
  assign tmp8453 = 1'b0;
  wire tmp8454;
  assign tmp8454 = (tmp8451 & tmp8452) | (tmp8451 & tmp8453) | (tmp8452 & tmp8453);
  wire tmp8455;
  assign tmp8455 = 1'b0;
  wire tmp8456;
  assign tmp8456 = 1'b0;
  wire tmp8457;
  assign tmp8457 = 1'b0;
  wire tmp8458;
  assign tmp8458 = (tmp8455 & tmp8456) | (tmp8455 & tmp8457) | (tmp8456 & tmp8457);
  wire tmp8459;
  assign tmp8459 = (tmp8450 & tmp8454) | (tmp8450 & tmp8458) | (tmp8454 & tmp8458);
  wire tmp8460;
  assign tmp8460 = (tmp8433 & tmp8446) | (tmp8433 & tmp8459) | (tmp8446 & tmp8459);
  wire tmp8461;
  assign tmp8461 = 1'b0;
  wire tmp8462;
  assign tmp8462 = 1'b0;
  wire tmp8463;
  assign tmp8463 = 1'b0;
  wire tmp8464;
  assign tmp8464 = (tmp8461 & tmp8462) | (tmp8461 & tmp8463) | (tmp8462 & tmp8463);
  wire tmp8465;
  assign tmp8465 = 1'b0;
  wire tmp8466;
  assign tmp8466 = 1'b0;
  wire tmp8467;
  assign tmp8467 = 1'b0;
  wire tmp8468;
  assign tmp8468 = (tmp8465 & tmp8466) | (tmp8465 & tmp8467) | (tmp8466 & tmp8467);
  wire tmp8469;
  assign tmp8469 = 1'b0;
  wire tmp8470;
  assign tmp8470 = 1'b0;
  wire tmp8471;
  assign tmp8471 = 1'b0;
  wire tmp8472;
  assign tmp8472 = (tmp8469 & tmp8470) | (tmp8469 & tmp8471) | (tmp8470 & tmp8471);
  wire tmp8473;
  assign tmp8473 = (tmp8464 & tmp8468) | (tmp8464 & tmp8472) | (tmp8468 & tmp8472);
  wire tmp8474;
  assign tmp8474 = 1'b0;
  wire tmp8475;
  assign tmp8475 = 1'b0;
  wire tmp8476;
  assign tmp8476 = 1'b0;
  wire tmp8477;
  assign tmp8477 = (tmp8474 & tmp8475) | (tmp8474 & tmp8476) | (tmp8475 & tmp8476);
  wire tmp8478;
  assign tmp8478 = 1'b0;
  wire tmp8479;
  assign tmp8479 = ~pi7;
  wire tmp8480;
  assign tmp8480 = 1'b0;
  wire tmp8481;
  assign tmp8481 = (tmp8478 & tmp8479) | (tmp8478 & tmp8480) | (tmp8479 & tmp8480);
  wire tmp8482;
  assign tmp8482 = 1'b0;
  wire tmp8483;
  assign tmp8483 = 1'b0;
  wire tmp8484;
  assign tmp8484 = 1'b0;
  wire tmp8485;
  assign tmp8485 = (tmp8482 & tmp8483) | (tmp8482 & tmp8484) | (tmp8483 & tmp8484);
  wire tmp8486;
  assign tmp8486 = (tmp8477 & tmp8481) | (tmp8477 & tmp8485) | (tmp8481 & tmp8485);
  wire tmp8487;
  assign tmp8487 = 1'b0;
  wire tmp8488;
  assign tmp8488 = 1'b0;
  wire tmp8489;
  assign tmp8489 = 1'b0;
  wire tmp8490;
  assign tmp8490 = (tmp8487 & tmp8488) | (tmp8487 & tmp8489) | (tmp8488 & tmp8489);
  wire tmp8491;
  assign tmp8491 = 1'b0;
  wire tmp8492;
  assign tmp8492 = 1'b0;
  wire tmp8493;
  assign tmp8493 = 1'b0;
  wire tmp8494;
  assign tmp8494 = (tmp8491 & tmp8492) | (tmp8491 & tmp8493) | (tmp8492 & tmp8493);
  wire tmp8495;
  assign tmp8495 = 1'b0;
  wire tmp8496;
  assign tmp8496 = 1'b0;
  wire tmp8497;
  assign tmp8497 = 1'b0;
  wire tmp8498;
  assign tmp8498 = (tmp8495 & tmp8496) | (tmp8495 & tmp8497) | (tmp8496 & tmp8497);
  wire tmp8499;
  assign tmp8499 = (tmp8490 & tmp8494) | (tmp8490 & tmp8498) | (tmp8494 & tmp8498);
  wire tmp8500;
  assign tmp8500 = (tmp8473 & tmp8486) | (tmp8473 & tmp8499) | (tmp8486 & tmp8499);
  wire tmp8501;
  assign tmp8501 = (tmp8420 & tmp8460) | (tmp8420 & tmp8500) | (tmp8460 & tmp8500);
  wire tmp8502;
  assign tmp8502 = 1'b0;
  wire tmp8503;
  assign tmp8503 = 1'b0;
  wire tmp8504;
  assign tmp8504 = 1'b0;
  wire tmp8505;
  assign tmp8505 = (tmp8502 & tmp8503) | (tmp8502 & tmp8504) | (tmp8503 & tmp8504);
  wire tmp8506;
  assign tmp8506 = 1'b0;
  wire tmp8507;
  assign tmp8507 = 1'b1;
  wire tmp8508;
  assign tmp8508 = 1'b0;
  wire tmp8509;
  assign tmp8509 = (tmp8506 & tmp8507) | (tmp8506 & tmp8508) | (tmp8507 & tmp8508);
  wire tmp8510;
  assign tmp8510 = 1'b0;
  wire tmp8511;
  assign tmp8511 = 1'b0;
  wire tmp8512;
  assign tmp8512 = 1'b0;
  wire tmp8513;
  assign tmp8513 = (tmp8510 & tmp8511) | (tmp8510 & tmp8512) | (tmp8511 & tmp8512);
  wire tmp8514;
  assign tmp8514 = (tmp8505 & tmp8509) | (tmp8505 & tmp8513) | (tmp8509 & tmp8513);
  wire tmp8515;
  assign tmp8515 = 1'b0;
  wire tmp8516;
  assign tmp8516 = 1'b1;
  wire tmp8517;
  assign tmp8517 = 1'b0;
  wire tmp8518;
  assign tmp8518 = (tmp8515 & tmp8516) | (tmp8515 & tmp8517) | (tmp8516 & tmp8517);
  wire tmp8519;
  assign tmp8519 = 1'b1;
  wire tmp8520;
  assign tmp8520 = ~pi6;
  wire tmp8521;
  assign tmp8521 = ~pi7;
  wire tmp8522;
  assign tmp8522 = (tmp8519 & tmp8520) | (tmp8519 & tmp8521) | (tmp8520 & tmp8521);
  wire tmp8523;
  assign tmp8523 = 1'b0;
  wire tmp8524;
  assign tmp8524 = ~pi7;
  wire tmp8525;
  assign tmp8525 = 1'b0;
  wire tmp8526;
  assign tmp8526 = (tmp8523 & tmp8524) | (tmp8523 & tmp8525) | (tmp8524 & tmp8525);
  wire tmp8527;
  assign tmp8527 = (tmp8518 & tmp8522) | (tmp8518 & tmp8526) | (tmp8522 & tmp8526);
  wire tmp8528;
  assign tmp8528 = 1'b0;
  wire tmp8529;
  assign tmp8529 = 1'b0;
  wire tmp8530;
  assign tmp8530 = 1'b0;
  wire tmp8531;
  assign tmp8531 = (tmp8528 & tmp8529) | (tmp8528 & tmp8530) | (tmp8529 & tmp8530);
  wire tmp8532;
  assign tmp8532 = 1'b0;
  wire tmp8533;
  assign tmp8533 = ~pi7;
  wire tmp8534;
  assign tmp8534 = 1'b0;
  wire tmp8535;
  assign tmp8535 = (tmp8532 & tmp8533) | (tmp8532 & tmp8534) | (tmp8533 & tmp8534);
  wire tmp8536;
  assign tmp8536 = 1'b0;
  wire tmp8537;
  assign tmp8537 = 1'b0;
  wire tmp8538;
  assign tmp8538 = 1'b0;
  wire tmp8539;
  assign tmp8539 = (tmp8536 & tmp8537) | (tmp8536 & tmp8538) | (tmp8537 & tmp8538);
  wire tmp8540;
  assign tmp8540 = (tmp8531 & tmp8535) | (tmp8531 & tmp8539) | (tmp8535 & tmp8539);
  wire tmp8541;
  assign tmp8541 = (tmp8514 & tmp8527) | (tmp8514 & tmp8540) | (tmp8527 & tmp8540);
  wire tmp8542;
  assign tmp8542 = 1'b0;
  wire tmp8543;
  assign tmp8543 = 1'b1;
  wire tmp8544;
  assign tmp8544 = 1'b0;
  wire tmp8545;
  assign tmp8545 = (tmp8542 & tmp8543) | (tmp8542 & tmp8544) | (tmp8543 & tmp8544);
  wire tmp8546;
  assign tmp8546 = 1'b1;
  wire tmp8547;
  assign tmp8547 = ~pi6;
  wire tmp8548;
  assign tmp8548 = ~pi7;
  wire tmp8549;
  assign tmp8549 = (tmp8546 & tmp8547) | (tmp8546 & tmp8548) | (tmp8547 & tmp8548);
  wire tmp8550;
  assign tmp8550 = 1'b0;
  wire tmp8551;
  assign tmp8551 = ~pi7;
  wire tmp8552;
  assign tmp8552 = 1'b0;
  wire tmp8553;
  assign tmp8553 = (tmp8550 & tmp8551) | (tmp8550 & tmp8552) | (tmp8551 & tmp8552);
  wire tmp8554;
  assign tmp8554 = (tmp8545 & tmp8549) | (tmp8545 & tmp8553) | (tmp8549 & tmp8553);
  wire tmp8555;
  assign tmp8555 = 1'b1;
  wire tmp8556;
  assign tmp8556 = ~pi6;
  wire tmp8557;
  assign tmp8557 = ~pi7;
  wire tmp8558;
  assign tmp8558 = (tmp8555 & tmp8556) | (tmp8555 & tmp8557) | (tmp8556 & tmp8557);
  wire tmp8559;
  assign tmp8559 = ~pi6;
  wire tmp8560;
  assign tmp8560 = 1'b1;
  wire tmp8561;
  assign tmp8561 = 1'b1;
  wire tmp8562;
  assign tmp8562 = (tmp8559 & tmp8560) | (tmp8559 & tmp8561) | (tmp8560 & tmp8561);
  wire tmp8563;
  assign tmp8563 = ~pi7;
  wire tmp8564;
  assign tmp8564 = 1'b1;
  wire tmp8565;
  assign tmp8565 = 1'b0;
  wire tmp8566;
  assign tmp8566 = (tmp8563 & tmp8564) | (tmp8563 & tmp8565) | (tmp8564 & tmp8565);
  wire tmp8567;
  assign tmp8567 = (tmp8558 & tmp8562) | (tmp8558 & tmp8566) | (tmp8562 & tmp8566);
  wire tmp8568;
  assign tmp8568 = 1'b0;
  wire tmp8569;
  assign tmp8569 = ~pi7;
  wire tmp8570;
  assign tmp8570 = 1'b0;
  wire tmp8571;
  assign tmp8571 = (tmp8568 & tmp8569) | (tmp8568 & tmp8570) | (tmp8569 & tmp8570);
  wire tmp8572;
  assign tmp8572 = ~pi7;
  wire tmp8573;
  assign tmp8573 = 1'b1;
  wire tmp8574;
  assign tmp8574 = 1'b0;
  wire tmp8575;
  assign tmp8575 = (tmp8572 & tmp8573) | (tmp8572 & tmp8574) | (tmp8573 & tmp8574);
  wire tmp8576;
  assign tmp8576 = 1'b0;
  wire tmp8577;
  assign tmp8577 = 1'b0;
  wire tmp8578;
  assign tmp8578 = 1'b0;
  wire tmp8579;
  assign tmp8579 = (tmp8576 & tmp8577) | (tmp8576 & tmp8578) | (tmp8577 & tmp8578);
  wire tmp8580;
  assign tmp8580 = (tmp8571 & tmp8575) | (tmp8571 & tmp8579) | (tmp8575 & tmp8579);
  wire tmp8581;
  assign tmp8581 = (tmp8554 & tmp8567) | (tmp8554 & tmp8580) | (tmp8567 & tmp8580);
  wire tmp8582;
  assign tmp8582 = 1'b0;
  wire tmp8583;
  assign tmp8583 = 1'b0;
  wire tmp8584;
  assign tmp8584 = 1'b0;
  wire tmp8585;
  assign tmp8585 = (tmp8582 & tmp8583) | (tmp8582 & tmp8584) | (tmp8583 & tmp8584);
  wire tmp8586;
  assign tmp8586 = 1'b0;
  wire tmp8587;
  assign tmp8587 = ~pi7;
  wire tmp8588;
  assign tmp8588 = 1'b0;
  wire tmp8589;
  assign tmp8589 = (tmp8586 & tmp8587) | (tmp8586 & tmp8588) | (tmp8587 & tmp8588);
  wire tmp8590;
  assign tmp8590 = 1'b0;
  wire tmp8591;
  assign tmp8591 = 1'b0;
  wire tmp8592;
  assign tmp8592 = 1'b0;
  wire tmp8593;
  assign tmp8593 = (tmp8590 & tmp8591) | (tmp8590 & tmp8592) | (tmp8591 & tmp8592);
  wire tmp8594;
  assign tmp8594 = (tmp8585 & tmp8589) | (tmp8585 & tmp8593) | (tmp8589 & tmp8593);
  wire tmp8595;
  assign tmp8595 = 1'b0;
  wire tmp8596;
  assign tmp8596 = ~pi7;
  wire tmp8597;
  assign tmp8597 = 1'b0;
  wire tmp8598;
  assign tmp8598 = (tmp8595 & tmp8596) | (tmp8595 & tmp8597) | (tmp8596 & tmp8597);
  wire tmp8599;
  assign tmp8599 = ~pi7;
  wire tmp8600;
  assign tmp8600 = 1'b1;
  wire tmp8601;
  assign tmp8601 = 1'b0;
  wire tmp8602;
  assign tmp8602 = (tmp8599 & tmp8600) | (tmp8599 & tmp8601) | (tmp8600 & tmp8601);
  wire tmp8603;
  assign tmp8603 = 1'b0;
  wire tmp8604;
  assign tmp8604 = 1'b0;
  wire tmp8605;
  assign tmp8605 = 1'b0;
  wire tmp8606;
  assign tmp8606 = (tmp8603 & tmp8604) | (tmp8603 & tmp8605) | (tmp8604 & tmp8605);
  wire tmp8607;
  assign tmp8607 = (tmp8598 & tmp8602) | (tmp8598 & tmp8606) | (tmp8602 & tmp8606);
  wire tmp8608;
  assign tmp8608 = 1'b0;
  wire tmp8609;
  assign tmp8609 = 1'b0;
  wire tmp8610;
  assign tmp8610 = 1'b0;
  wire tmp8611;
  assign tmp8611 = (tmp8608 & tmp8609) | (tmp8608 & tmp8610) | (tmp8609 & tmp8610);
  wire tmp8612;
  assign tmp8612 = 1'b0;
  wire tmp8613;
  assign tmp8613 = 1'b0;
  wire tmp8614;
  assign tmp8614 = 1'b0;
  wire tmp8615;
  assign tmp8615 = (tmp8612 & tmp8613) | (tmp8612 & tmp8614) | (tmp8613 & tmp8614);
  wire tmp8616;
  assign tmp8616 = 1'b0;
  wire tmp8617;
  assign tmp8617 = 1'b0;
  wire tmp8618;
  assign tmp8618 = 1'b0;
  wire tmp8619;
  assign tmp8619 = (tmp8616 & tmp8617) | (tmp8616 & tmp8618) | (tmp8617 & tmp8618);
  wire tmp8620;
  assign tmp8620 = (tmp8611 & tmp8615) | (tmp8611 & tmp8619) | (tmp8615 & tmp8619);
  wire tmp8621;
  assign tmp8621 = (tmp8594 & tmp8607) | (tmp8594 & tmp8620) | (tmp8607 & tmp8620);
  wire tmp8622;
  assign tmp8622 = (tmp8541 & tmp8581) | (tmp8541 & tmp8621) | (tmp8581 & tmp8621);
  wire tmp8623;
  assign tmp8623 = 1'b0;
  wire tmp8624;
  assign tmp8624 = 1'b0;
  wire tmp8625;
  assign tmp8625 = 1'b0;
  wire tmp8626;
  assign tmp8626 = (tmp8623 & tmp8624) | (tmp8623 & tmp8625) | (tmp8624 & tmp8625);
  wire tmp8627;
  assign tmp8627 = 1'b0;
  wire tmp8628;
  assign tmp8628 = 1'b0;
  wire tmp8629;
  assign tmp8629 = 1'b0;
  wire tmp8630;
  assign tmp8630 = (tmp8627 & tmp8628) | (tmp8627 & tmp8629) | (tmp8628 & tmp8629);
  wire tmp8631;
  assign tmp8631 = 1'b0;
  wire tmp8632;
  assign tmp8632 = 1'b0;
  wire tmp8633;
  assign tmp8633 = 1'b0;
  wire tmp8634;
  assign tmp8634 = (tmp8631 & tmp8632) | (tmp8631 & tmp8633) | (tmp8632 & tmp8633);
  wire tmp8635;
  assign tmp8635 = (tmp8626 & tmp8630) | (tmp8626 & tmp8634) | (tmp8630 & tmp8634);
  wire tmp8636;
  assign tmp8636 = 1'b0;
  wire tmp8637;
  assign tmp8637 = 1'b0;
  wire tmp8638;
  assign tmp8638 = 1'b0;
  wire tmp8639;
  assign tmp8639 = (tmp8636 & tmp8637) | (tmp8636 & tmp8638) | (tmp8637 & tmp8638);
  wire tmp8640;
  assign tmp8640 = 1'b0;
  wire tmp8641;
  assign tmp8641 = ~pi7;
  wire tmp8642;
  assign tmp8642 = 1'b0;
  wire tmp8643;
  assign tmp8643 = (tmp8640 & tmp8641) | (tmp8640 & tmp8642) | (tmp8641 & tmp8642);
  wire tmp8644;
  assign tmp8644 = 1'b0;
  wire tmp8645;
  assign tmp8645 = 1'b0;
  wire tmp8646;
  assign tmp8646 = 1'b0;
  wire tmp8647;
  assign tmp8647 = (tmp8644 & tmp8645) | (tmp8644 & tmp8646) | (tmp8645 & tmp8646);
  wire tmp8648;
  assign tmp8648 = (tmp8639 & tmp8643) | (tmp8639 & tmp8647) | (tmp8643 & tmp8647);
  wire tmp8649;
  assign tmp8649 = 1'b0;
  wire tmp8650;
  assign tmp8650 = 1'b0;
  wire tmp8651;
  assign tmp8651 = 1'b0;
  wire tmp8652;
  assign tmp8652 = (tmp8649 & tmp8650) | (tmp8649 & tmp8651) | (tmp8650 & tmp8651);
  wire tmp8653;
  assign tmp8653 = 1'b0;
  wire tmp8654;
  assign tmp8654 = 1'b0;
  wire tmp8655;
  assign tmp8655 = 1'b0;
  wire tmp8656;
  assign tmp8656 = (tmp8653 & tmp8654) | (tmp8653 & tmp8655) | (tmp8654 & tmp8655);
  wire tmp8657;
  assign tmp8657 = 1'b0;
  wire tmp8658;
  assign tmp8658 = 1'b0;
  wire tmp8659;
  assign tmp8659 = 1'b0;
  wire tmp8660;
  assign tmp8660 = (tmp8657 & tmp8658) | (tmp8657 & tmp8659) | (tmp8658 & tmp8659);
  wire tmp8661;
  assign tmp8661 = (tmp8652 & tmp8656) | (tmp8652 & tmp8660) | (tmp8656 & tmp8660);
  wire tmp8662;
  assign tmp8662 = (tmp8635 & tmp8648) | (tmp8635 & tmp8661) | (tmp8648 & tmp8661);
  wire tmp8663;
  assign tmp8663 = 1'b0;
  wire tmp8664;
  assign tmp8664 = 1'b0;
  wire tmp8665;
  assign tmp8665 = 1'b0;
  wire tmp8666;
  assign tmp8666 = (tmp8663 & tmp8664) | (tmp8663 & tmp8665) | (tmp8664 & tmp8665);
  wire tmp8667;
  assign tmp8667 = 1'b0;
  wire tmp8668;
  assign tmp8668 = ~pi7;
  wire tmp8669;
  assign tmp8669 = 1'b0;
  wire tmp8670;
  assign tmp8670 = (tmp8667 & tmp8668) | (tmp8667 & tmp8669) | (tmp8668 & tmp8669);
  wire tmp8671;
  assign tmp8671 = 1'b0;
  wire tmp8672;
  assign tmp8672 = 1'b0;
  wire tmp8673;
  assign tmp8673 = 1'b0;
  wire tmp8674;
  assign tmp8674 = (tmp8671 & tmp8672) | (tmp8671 & tmp8673) | (tmp8672 & tmp8673);
  wire tmp8675;
  assign tmp8675 = (tmp8666 & tmp8670) | (tmp8666 & tmp8674) | (tmp8670 & tmp8674);
  wire tmp8676;
  assign tmp8676 = 1'b0;
  wire tmp8677;
  assign tmp8677 = ~pi7;
  wire tmp8678;
  assign tmp8678 = 1'b0;
  wire tmp8679;
  assign tmp8679 = (tmp8676 & tmp8677) | (tmp8676 & tmp8678) | (tmp8677 & tmp8678);
  wire tmp8680;
  assign tmp8680 = ~pi7;
  wire tmp8681;
  assign tmp8681 = 1'b1;
  wire tmp8682;
  assign tmp8682 = 1'b0;
  wire tmp8683;
  assign tmp8683 = (tmp8680 & tmp8681) | (tmp8680 & tmp8682) | (tmp8681 & tmp8682);
  wire tmp8684;
  assign tmp8684 = 1'b0;
  wire tmp8685;
  assign tmp8685 = 1'b0;
  wire tmp8686;
  assign tmp8686 = 1'b0;
  wire tmp8687;
  assign tmp8687 = (tmp8684 & tmp8685) | (tmp8684 & tmp8686) | (tmp8685 & tmp8686);
  wire tmp8688;
  assign tmp8688 = (tmp8679 & tmp8683) | (tmp8679 & tmp8687) | (tmp8683 & tmp8687);
  wire tmp8689;
  assign tmp8689 = 1'b0;
  wire tmp8690;
  assign tmp8690 = 1'b0;
  wire tmp8691;
  assign tmp8691 = 1'b0;
  wire tmp8692;
  assign tmp8692 = (tmp8689 & tmp8690) | (tmp8689 & tmp8691) | (tmp8690 & tmp8691);
  wire tmp8693;
  assign tmp8693 = 1'b0;
  wire tmp8694;
  assign tmp8694 = 1'b0;
  wire tmp8695;
  assign tmp8695 = 1'b0;
  wire tmp8696;
  assign tmp8696 = (tmp8693 & tmp8694) | (tmp8693 & tmp8695) | (tmp8694 & tmp8695);
  wire tmp8697;
  assign tmp8697 = 1'b0;
  wire tmp8698;
  assign tmp8698 = 1'b0;
  wire tmp8699;
  assign tmp8699 = 1'b0;
  wire tmp8700;
  assign tmp8700 = (tmp8697 & tmp8698) | (tmp8697 & tmp8699) | (tmp8698 & tmp8699);
  wire tmp8701;
  assign tmp8701 = (tmp8692 & tmp8696) | (tmp8692 & tmp8700) | (tmp8696 & tmp8700);
  wire tmp8702;
  assign tmp8702 = (tmp8675 & tmp8688) | (tmp8675 & tmp8701) | (tmp8688 & tmp8701);
  wire tmp8703;
  assign tmp8703 = 1'b0;
  wire tmp8704;
  assign tmp8704 = 1'b0;
  wire tmp8705;
  assign tmp8705 = 1'b0;
  wire tmp8706;
  assign tmp8706 = (tmp8703 & tmp8704) | (tmp8703 & tmp8705) | (tmp8704 & tmp8705);
  wire tmp8707;
  assign tmp8707 = 1'b0;
  wire tmp8708;
  assign tmp8708 = 1'b0;
  wire tmp8709;
  assign tmp8709 = 1'b0;
  wire tmp8710;
  assign tmp8710 = (tmp8707 & tmp8708) | (tmp8707 & tmp8709) | (tmp8708 & tmp8709);
  wire tmp8711;
  assign tmp8711 = 1'b0;
  wire tmp8712;
  assign tmp8712 = 1'b0;
  wire tmp8713;
  assign tmp8713 = 1'b0;
  wire tmp8714;
  assign tmp8714 = (tmp8711 & tmp8712) | (tmp8711 & tmp8713) | (tmp8712 & tmp8713);
  wire tmp8715;
  assign tmp8715 = (tmp8706 & tmp8710) | (tmp8706 & tmp8714) | (tmp8710 & tmp8714);
  wire tmp8716;
  assign tmp8716 = 1'b0;
  wire tmp8717;
  assign tmp8717 = 1'b0;
  wire tmp8718;
  assign tmp8718 = 1'b0;
  wire tmp8719;
  assign tmp8719 = (tmp8716 & tmp8717) | (tmp8716 & tmp8718) | (tmp8717 & tmp8718);
  wire tmp8720;
  assign tmp8720 = 1'b0;
  wire tmp8721;
  assign tmp8721 = 1'b0;
  wire tmp8722;
  assign tmp8722 = 1'b0;
  wire tmp8723;
  assign tmp8723 = (tmp8720 & tmp8721) | (tmp8720 & tmp8722) | (tmp8721 & tmp8722);
  wire tmp8724;
  assign tmp8724 = 1'b0;
  wire tmp8725;
  assign tmp8725 = 1'b0;
  wire tmp8726;
  assign tmp8726 = 1'b0;
  wire tmp8727;
  assign tmp8727 = (tmp8724 & tmp8725) | (tmp8724 & tmp8726) | (tmp8725 & tmp8726);
  wire tmp8728;
  assign tmp8728 = (tmp8719 & tmp8723) | (tmp8719 & tmp8727) | (tmp8723 & tmp8727);
  wire tmp8729;
  assign tmp8729 = 1'b0;
  wire tmp8730;
  assign tmp8730 = 1'b0;
  wire tmp8731;
  assign tmp8731 = 1'b0;
  wire tmp8732;
  assign tmp8732 = (tmp8729 & tmp8730) | (tmp8729 & tmp8731) | (tmp8730 & tmp8731);
  wire tmp8733;
  assign tmp8733 = 1'b0;
  wire tmp8734;
  assign tmp8734 = 1'b0;
  wire tmp8735;
  assign tmp8735 = 1'b0;
  wire tmp8736;
  assign tmp8736 = (tmp8733 & tmp8734) | (tmp8733 & tmp8735) | (tmp8734 & tmp8735);
  wire tmp8737;
  assign tmp8737 = 1'b0;
  wire tmp8738;
  assign tmp8738 = 1'b0;
  wire tmp8739;
  assign tmp8739 = 1'b0;
  wire tmp8740;
  assign tmp8740 = (tmp8737 & tmp8738) | (tmp8737 & tmp8739) | (tmp8738 & tmp8739);
  wire tmp8741;
  assign tmp8741 = (tmp8732 & tmp8736) | (tmp8732 & tmp8740) | (tmp8736 & tmp8740);
  wire tmp8742;
  assign tmp8742 = (tmp8715 & tmp8728) | (tmp8715 & tmp8741) | (tmp8728 & tmp8741);
  wire tmp8743;
  assign tmp8743 = (tmp8662 & tmp8702) | (tmp8662 & tmp8742) | (tmp8702 & tmp8742);
  wire tmp8744;
  assign tmp8744 = (tmp8501 & tmp8622) | (tmp8501 & tmp8743) | (tmp8622 & tmp8743);
  wire tmp8745;
  assign tmp8745 = (tmp8016 & tmp8380) | (tmp8016 & tmp8744) | (tmp8380 & tmp8744);
  wire tmp8746;
  assign tmp8746 = 1'b0;
  wire tmp8747;
  assign tmp8747 = 1'b0;
  wire tmp8748;
  assign tmp8748 = 1'b0;
  wire tmp8749;
  assign tmp8749 = (tmp8746 & tmp8747) | (tmp8746 & tmp8748) | (tmp8747 & tmp8748);
  wire tmp8750;
  assign tmp8750 = 1'b0;
  wire tmp8751;
  assign tmp8751 = 1'b0;
  wire tmp8752;
  assign tmp8752 = 1'b0;
  wire tmp8753;
  assign tmp8753 = (tmp8750 & tmp8751) | (tmp8750 & tmp8752) | (tmp8751 & tmp8752);
  wire tmp8754;
  assign tmp8754 = 1'b0;
  wire tmp8755;
  assign tmp8755 = 1'b0;
  wire tmp8756;
  assign tmp8756 = 1'b0;
  wire tmp8757;
  assign tmp8757 = (tmp8754 & tmp8755) | (tmp8754 & tmp8756) | (tmp8755 & tmp8756);
  wire tmp8758;
  assign tmp8758 = (tmp8749 & tmp8753) | (tmp8749 & tmp8757) | (tmp8753 & tmp8757);
  wire tmp8759;
  assign tmp8759 = 1'b0;
  wire tmp8760;
  assign tmp8760 = 1'b0;
  wire tmp8761;
  assign tmp8761 = 1'b0;
  wire tmp8762;
  assign tmp8762 = (tmp8759 & tmp8760) | (tmp8759 & tmp8761) | (tmp8760 & tmp8761);
  wire tmp8763;
  assign tmp8763 = 1'b0;
  wire tmp8764;
  assign tmp8764 = 1'b0;
  wire tmp8765;
  assign tmp8765 = 1'b0;
  wire tmp8766;
  assign tmp8766 = (tmp8763 & tmp8764) | (tmp8763 & tmp8765) | (tmp8764 & tmp8765);
  wire tmp8767;
  assign tmp8767 = 1'b0;
  wire tmp8768;
  assign tmp8768 = 1'b0;
  wire tmp8769;
  assign tmp8769 = 1'b0;
  wire tmp8770;
  assign tmp8770 = (tmp8767 & tmp8768) | (tmp8767 & tmp8769) | (tmp8768 & tmp8769);
  wire tmp8771;
  assign tmp8771 = (tmp8762 & tmp8766) | (tmp8762 & tmp8770) | (tmp8766 & tmp8770);
  wire tmp8772;
  assign tmp8772 = 1'b0;
  wire tmp8773;
  assign tmp8773 = 1'b0;
  wire tmp8774;
  assign tmp8774 = 1'b0;
  wire tmp8775;
  assign tmp8775 = (tmp8772 & tmp8773) | (tmp8772 & tmp8774) | (tmp8773 & tmp8774);
  wire tmp8776;
  assign tmp8776 = 1'b0;
  wire tmp8777;
  assign tmp8777 = 1'b0;
  wire tmp8778;
  assign tmp8778 = 1'b0;
  wire tmp8779;
  assign tmp8779 = (tmp8776 & tmp8777) | (tmp8776 & tmp8778) | (tmp8777 & tmp8778);
  wire tmp8780;
  assign tmp8780 = 1'b0;
  wire tmp8781;
  assign tmp8781 = 1'b0;
  wire tmp8782;
  assign tmp8782 = 1'b0;
  wire tmp8783;
  assign tmp8783 = (tmp8780 & tmp8781) | (tmp8780 & tmp8782) | (tmp8781 & tmp8782);
  wire tmp8784;
  assign tmp8784 = (tmp8775 & tmp8779) | (tmp8775 & tmp8783) | (tmp8779 & tmp8783);
  wire tmp8785;
  assign tmp8785 = (tmp8758 & tmp8771) | (tmp8758 & tmp8784) | (tmp8771 & tmp8784);
  wire tmp8786;
  assign tmp8786 = 1'b0;
  wire tmp8787;
  assign tmp8787 = 1'b0;
  wire tmp8788;
  assign tmp8788 = 1'b0;
  wire tmp8789;
  assign tmp8789 = (tmp8786 & tmp8787) | (tmp8786 & tmp8788) | (tmp8787 & tmp8788);
  wire tmp8790;
  assign tmp8790 = 1'b0;
  wire tmp8791;
  assign tmp8791 = 1'b0;
  wire tmp8792;
  assign tmp8792 = 1'b0;
  wire tmp8793;
  assign tmp8793 = (tmp8790 & tmp8791) | (tmp8790 & tmp8792) | (tmp8791 & tmp8792);
  wire tmp8794;
  assign tmp8794 = 1'b0;
  wire tmp8795;
  assign tmp8795 = 1'b0;
  wire tmp8796;
  assign tmp8796 = 1'b0;
  wire tmp8797;
  assign tmp8797 = (tmp8794 & tmp8795) | (tmp8794 & tmp8796) | (tmp8795 & tmp8796);
  wire tmp8798;
  assign tmp8798 = (tmp8789 & tmp8793) | (tmp8789 & tmp8797) | (tmp8793 & tmp8797);
  wire tmp8799;
  assign tmp8799 = 1'b0;
  wire tmp8800;
  assign tmp8800 = 1'b0;
  wire tmp8801;
  assign tmp8801 = 1'b0;
  wire tmp8802;
  assign tmp8802 = (tmp8799 & tmp8800) | (tmp8799 & tmp8801) | (tmp8800 & tmp8801);
  wire tmp8803;
  assign tmp8803 = 1'b0;
  wire tmp8804;
  assign tmp8804 = 1'b1;
  wire tmp8805;
  assign tmp8805 = 1'b0;
  wire tmp8806;
  assign tmp8806 = (tmp8803 & tmp8804) | (tmp8803 & tmp8805) | (tmp8804 & tmp8805);
  wire tmp8807;
  assign tmp8807 = 1'b0;
  wire tmp8808;
  assign tmp8808 = 1'b0;
  wire tmp8809;
  assign tmp8809 = 1'b0;
  wire tmp8810;
  assign tmp8810 = (tmp8807 & tmp8808) | (tmp8807 & tmp8809) | (tmp8808 & tmp8809);
  wire tmp8811;
  assign tmp8811 = (tmp8802 & tmp8806) | (tmp8802 & tmp8810) | (tmp8806 & tmp8810);
  wire tmp8812;
  assign tmp8812 = 1'b0;
  wire tmp8813;
  assign tmp8813 = 1'b0;
  wire tmp8814;
  assign tmp8814 = 1'b0;
  wire tmp8815;
  assign tmp8815 = (tmp8812 & tmp8813) | (tmp8812 & tmp8814) | (tmp8813 & tmp8814);
  wire tmp8816;
  assign tmp8816 = 1'b0;
  wire tmp8817;
  assign tmp8817 = 1'b0;
  wire tmp8818;
  assign tmp8818 = 1'b0;
  wire tmp8819;
  assign tmp8819 = (tmp8816 & tmp8817) | (tmp8816 & tmp8818) | (tmp8817 & tmp8818);
  wire tmp8820;
  assign tmp8820 = 1'b0;
  wire tmp8821;
  assign tmp8821 = 1'b0;
  wire tmp8822;
  assign tmp8822 = 1'b0;
  wire tmp8823;
  assign tmp8823 = (tmp8820 & tmp8821) | (tmp8820 & tmp8822) | (tmp8821 & tmp8822);
  wire tmp8824;
  assign tmp8824 = (tmp8815 & tmp8819) | (tmp8815 & tmp8823) | (tmp8819 & tmp8823);
  wire tmp8825;
  assign tmp8825 = (tmp8798 & tmp8811) | (tmp8798 & tmp8824) | (tmp8811 & tmp8824);
  wire tmp8826;
  assign tmp8826 = 1'b0;
  wire tmp8827;
  assign tmp8827 = 1'b0;
  wire tmp8828;
  assign tmp8828 = 1'b0;
  wire tmp8829;
  assign tmp8829 = (tmp8826 & tmp8827) | (tmp8826 & tmp8828) | (tmp8827 & tmp8828);
  wire tmp8830;
  assign tmp8830 = 1'b0;
  wire tmp8831;
  assign tmp8831 = 1'b0;
  wire tmp8832;
  assign tmp8832 = 1'b0;
  wire tmp8833;
  assign tmp8833 = (tmp8830 & tmp8831) | (tmp8830 & tmp8832) | (tmp8831 & tmp8832);
  wire tmp8834;
  assign tmp8834 = 1'b0;
  wire tmp8835;
  assign tmp8835 = 1'b0;
  wire tmp8836;
  assign tmp8836 = 1'b0;
  wire tmp8837;
  assign tmp8837 = (tmp8834 & tmp8835) | (tmp8834 & tmp8836) | (tmp8835 & tmp8836);
  wire tmp8838;
  assign tmp8838 = (tmp8829 & tmp8833) | (tmp8829 & tmp8837) | (tmp8833 & tmp8837);
  wire tmp8839;
  assign tmp8839 = 1'b0;
  wire tmp8840;
  assign tmp8840 = 1'b0;
  wire tmp8841;
  assign tmp8841 = 1'b0;
  wire tmp8842;
  assign tmp8842 = (tmp8839 & tmp8840) | (tmp8839 & tmp8841) | (tmp8840 & tmp8841);
  wire tmp8843;
  assign tmp8843 = 1'b0;
  wire tmp8844;
  assign tmp8844 = 1'b0;
  wire tmp8845;
  assign tmp8845 = 1'b0;
  wire tmp8846;
  assign tmp8846 = (tmp8843 & tmp8844) | (tmp8843 & tmp8845) | (tmp8844 & tmp8845);
  wire tmp8847;
  assign tmp8847 = 1'b0;
  wire tmp8848;
  assign tmp8848 = 1'b0;
  wire tmp8849;
  assign tmp8849 = 1'b0;
  wire tmp8850;
  assign tmp8850 = (tmp8847 & tmp8848) | (tmp8847 & tmp8849) | (tmp8848 & tmp8849);
  wire tmp8851;
  assign tmp8851 = (tmp8842 & tmp8846) | (tmp8842 & tmp8850) | (tmp8846 & tmp8850);
  wire tmp8852;
  assign tmp8852 = 1'b0;
  wire tmp8853;
  assign tmp8853 = 1'b0;
  wire tmp8854;
  assign tmp8854 = 1'b0;
  wire tmp8855;
  assign tmp8855 = (tmp8852 & tmp8853) | (tmp8852 & tmp8854) | (tmp8853 & tmp8854);
  wire tmp8856;
  assign tmp8856 = 1'b0;
  wire tmp8857;
  assign tmp8857 = 1'b0;
  wire tmp8858;
  assign tmp8858 = 1'b0;
  wire tmp8859;
  assign tmp8859 = (tmp8856 & tmp8857) | (tmp8856 & tmp8858) | (tmp8857 & tmp8858);
  wire tmp8860;
  assign tmp8860 = 1'b0;
  wire tmp8861;
  assign tmp8861 = 1'b0;
  wire tmp8862;
  assign tmp8862 = 1'b0;
  wire tmp8863;
  assign tmp8863 = (tmp8860 & tmp8861) | (tmp8860 & tmp8862) | (tmp8861 & tmp8862);
  wire tmp8864;
  assign tmp8864 = (tmp8855 & tmp8859) | (tmp8855 & tmp8863) | (tmp8859 & tmp8863);
  wire tmp8865;
  assign tmp8865 = (tmp8838 & tmp8851) | (tmp8838 & tmp8864) | (tmp8851 & tmp8864);
  wire tmp8866;
  assign tmp8866 = (tmp8785 & tmp8825) | (tmp8785 & tmp8865) | (tmp8825 & tmp8865);
  wire tmp8867;
  assign tmp8867 = 1'b0;
  wire tmp8868;
  assign tmp8868 = 1'b0;
  wire tmp8869;
  assign tmp8869 = 1'b0;
  wire tmp8870;
  assign tmp8870 = (tmp8867 & tmp8868) | (tmp8867 & tmp8869) | (tmp8868 & tmp8869);
  wire tmp8871;
  assign tmp8871 = 1'b0;
  wire tmp8872;
  assign tmp8872 = 1'b0;
  wire tmp8873;
  assign tmp8873 = 1'b0;
  wire tmp8874;
  assign tmp8874 = (tmp8871 & tmp8872) | (tmp8871 & tmp8873) | (tmp8872 & tmp8873);
  wire tmp8875;
  assign tmp8875 = 1'b0;
  wire tmp8876;
  assign tmp8876 = 1'b0;
  wire tmp8877;
  assign tmp8877 = 1'b0;
  wire tmp8878;
  assign tmp8878 = (tmp8875 & tmp8876) | (tmp8875 & tmp8877) | (tmp8876 & tmp8877);
  wire tmp8879;
  assign tmp8879 = (tmp8870 & tmp8874) | (tmp8870 & tmp8878) | (tmp8874 & tmp8878);
  wire tmp8880;
  assign tmp8880 = 1'b0;
  wire tmp8881;
  assign tmp8881 = 1'b0;
  wire tmp8882;
  assign tmp8882 = 1'b0;
  wire tmp8883;
  assign tmp8883 = (tmp8880 & tmp8881) | (tmp8880 & tmp8882) | (tmp8881 & tmp8882);
  wire tmp8884;
  assign tmp8884 = 1'b0;
  wire tmp8885;
  assign tmp8885 = 1'b1;
  wire tmp8886;
  assign tmp8886 = 1'b0;
  wire tmp8887;
  assign tmp8887 = (tmp8884 & tmp8885) | (tmp8884 & tmp8886) | (tmp8885 & tmp8886);
  wire tmp8888;
  assign tmp8888 = 1'b0;
  wire tmp8889;
  assign tmp8889 = 1'b0;
  wire tmp8890;
  assign tmp8890 = 1'b0;
  wire tmp8891;
  assign tmp8891 = (tmp8888 & tmp8889) | (tmp8888 & tmp8890) | (tmp8889 & tmp8890);
  wire tmp8892;
  assign tmp8892 = (tmp8883 & tmp8887) | (tmp8883 & tmp8891) | (tmp8887 & tmp8891);
  wire tmp8893;
  assign tmp8893 = 1'b0;
  wire tmp8894;
  assign tmp8894 = 1'b0;
  wire tmp8895;
  assign tmp8895 = 1'b0;
  wire tmp8896;
  assign tmp8896 = (tmp8893 & tmp8894) | (tmp8893 & tmp8895) | (tmp8894 & tmp8895);
  wire tmp8897;
  assign tmp8897 = 1'b0;
  wire tmp8898;
  assign tmp8898 = 1'b0;
  wire tmp8899;
  assign tmp8899 = 1'b0;
  wire tmp8900;
  assign tmp8900 = (tmp8897 & tmp8898) | (tmp8897 & tmp8899) | (tmp8898 & tmp8899);
  wire tmp8901;
  assign tmp8901 = 1'b0;
  wire tmp8902;
  assign tmp8902 = 1'b0;
  wire tmp8903;
  assign tmp8903 = 1'b0;
  wire tmp8904;
  assign tmp8904 = (tmp8901 & tmp8902) | (tmp8901 & tmp8903) | (tmp8902 & tmp8903);
  wire tmp8905;
  assign tmp8905 = (tmp8896 & tmp8900) | (tmp8896 & tmp8904) | (tmp8900 & tmp8904);
  wire tmp8906;
  assign tmp8906 = (tmp8879 & tmp8892) | (tmp8879 & tmp8905) | (tmp8892 & tmp8905);
  wire tmp8907;
  assign tmp8907 = 1'b0;
  wire tmp8908;
  assign tmp8908 = 1'b0;
  wire tmp8909;
  assign tmp8909 = 1'b0;
  wire tmp8910;
  assign tmp8910 = (tmp8907 & tmp8908) | (tmp8907 & tmp8909) | (tmp8908 & tmp8909);
  wire tmp8911;
  assign tmp8911 = 1'b0;
  wire tmp8912;
  assign tmp8912 = 1'b1;
  wire tmp8913;
  assign tmp8913 = 1'b0;
  wire tmp8914;
  assign tmp8914 = (tmp8911 & tmp8912) | (tmp8911 & tmp8913) | (tmp8912 & tmp8913);
  wire tmp8915;
  assign tmp8915 = 1'b0;
  wire tmp8916;
  assign tmp8916 = 1'b0;
  wire tmp8917;
  assign tmp8917 = 1'b0;
  wire tmp8918;
  assign tmp8918 = (tmp8915 & tmp8916) | (tmp8915 & tmp8917) | (tmp8916 & tmp8917);
  wire tmp8919;
  assign tmp8919 = (tmp8910 & tmp8914) | (tmp8910 & tmp8918) | (tmp8914 & tmp8918);
  wire tmp8920;
  assign tmp8920 = 1'b0;
  wire tmp8921;
  assign tmp8921 = 1'b1;
  wire tmp8922;
  assign tmp8922 = 1'b0;
  wire tmp8923;
  assign tmp8923 = (tmp8920 & tmp8921) | (tmp8920 & tmp8922) | (tmp8921 & tmp8922);
  wire tmp8924;
  assign tmp8924 = 1'b1;
  wire tmp8925;
  assign tmp8925 = ~pi6;
  wire tmp8926;
  assign tmp8926 = ~pi7;
  wire tmp8927;
  assign tmp8927 = (tmp8924 & tmp8925) | (tmp8924 & tmp8926) | (tmp8925 & tmp8926);
  wire tmp8928;
  assign tmp8928 = 1'b0;
  wire tmp8929;
  assign tmp8929 = ~pi7;
  wire tmp8930;
  assign tmp8930 = 1'b0;
  wire tmp8931;
  assign tmp8931 = (tmp8928 & tmp8929) | (tmp8928 & tmp8930) | (tmp8929 & tmp8930);
  wire tmp8932;
  assign tmp8932 = (tmp8923 & tmp8927) | (tmp8923 & tmp8931) | (tmp8927 & tmp8931);
  wire tmp8933;
  assign tmp8933 = 1'b0;
  wire tmp8934;
  assign tmp8934 = 1'b0;
  wire tmp8935;
  assign tmp8935 = 1'b0;
  wire tmp8936;
  assign tmp8936 = (tmp8933 & tmp8934) | (tmp8933 & tmp8935) | (tmp8934 & tmp8935);
  wire tmp8937;
  assign tmp8937 = 1'b0;
  wire tmp8938;
  assign tmp8938 = ~pi7;
  wire tmp8939;
  assign tmp8939 = 1'b0;
  wire tmp8940;
  assign tmp8940 = (tmp8937 & tmp8938) | (tmp8937 & tmp8939) | (tmp8938 & tmp8939);
  wire tmp8941;
  assign tmp8941 = 1'b0;
  wire tmp8942;
  assign tmp8942 = 1'b0;
  wire tmp8943;
  assign tmp8943 = 1'b0;
  wire tmp8944;
  assign tmp8944 = (tmp8941 & tmp8942) | (tmp8941 & tmp8943) | (tmp8942 & tmp8943);
  wire tmp8945;
  assign tmp8945 = (tmp8936 & tmp8940) | (tmp8936 & tmp8944) | (tmp8940 & tmp8944);
  wire tmp8946;
  assign tmp8946 = (tmp8919 & tmp8932) | (tmp8919 & tmp8945) | (tmp8932 & tmp8945);
  wire tmp8947;
  assign tmp8947 = 1'b0;
  wire tmp8948;
  assign tmp8948 = 1'b0;
  wire tmp8949;
  assign tmp8949 = 1'b0;
  wire tmp8950;
  assign tmp8950 = (tmp8947 & tmp8948) | (tmp8947 & tmp8949) | (tmp8948 & tmp8949);
  wire tmp8951;
  assign tmp8951 = 1'b0;
  wire tmp8952;
  assign tmp8952 = 1'b0;
  wire tmp8953;
  assign tmp8953 = 1'b0;
  wire tmp8954;
  assign tmp8954 = (tmp8951 & tmp8952) | (tmp8951 & tmp8953) | (tmp8952 & tmp8953);
  wire tmp8955;
  assign tmp8955 = 1'b0;
  wire tmp8956;
  assign tmp8956 = 1'b0;
  wire tmp8957;
  assign tmp8957 = 1'b0;
  wire tmp8958;
  assign tmp8958 = (tmp8955 & tmp8956) | (tmp8955 & tmp8957) | (tmp8956 & tmp8957);
  wire tmp8959;
  assign tmp8959 = (tmp8950 & tmp8954) | (tmp8950 & tmp8958) | (tmp8954 & tmp8958);
  wire tmp8960;
  assign tmp8960 = 1'b0;
  wire tmp8961;
  assign tmp8961 = 1'b0;
  wire tmp8962;
  assign tmp8962 = 1'b0;
  wire tmp8963;
  assign tmp8963 = (tmp8960 & tmp8961) | (tmp8960 & tmp8962) | (tmp8961 & tmp8962);
  wire tmp8964;
  assign tmp8964 = 1'b0;
  wire tmp8965;
  assign tmp8965 = ~pi7;
  wire tmp8966;
  assign tmp8966 = 1'b0;
  wire tmp8967;
  assign tmp8967 = (tmp8964 & tmp8965) | (tmp8964 & tmp8966) | (tmp8965 & tmp8966);
  wire tmp8968;
  assign tmp8968 = 1'b0;
  wire tmp8969;
  assign tmp8969 = 1'b0;
  wire tmp8970;
  assign tmp8970 = 1'b0;
  wire tmp8971;
  assign tmp8971 = (tmp8968 & tmp8969) | (tmp8968 & tmp8970) | (tmp8969 & tmp8970);
  wire tmp8972;
  assign tmp8972 = (tmp8963 & tmp8967) | (tmp8963 & tmp8971) | (tmp8967 & tmp8971);
  wire tmp8973;
  assign tmp8973 = 1'b0;
  wire tmp8974;
  assign tmp8974 = 1'b0;
  wire tmp8975;
  assign tmp8975 = 1'b0;
  wire tmp8976;
  assign tmp8976 = (tmp8973 & tmp8974) | (tmp8973 & tmp8975) | (tmp8974 & tmp8975);
  wire tmp8977;
  assign tmp8977 = 1'b0;
  wire tmp8978;
  assign tmp8978 = 1'b0;
  wire tmp8979;
  assign tmp8979 = 1'b0;
  wire tmp8980;
  assign tmp8980 = (tmp8977 & tmp8978) | (tmp8977 & tmp8979) | (tmp8978 & tmp8979);
  wire tmp8981;
  assign tmp8981 = 1'b0;
  wire tmp8982;
  assign tmp8982 = 1'b0;
  wire tmp8983;
  assign tmp8983 = 1'b0;
  wire tmp8984;
  assign tmp8984 = (tmp8981 & tmp8982) | (tmp8981 & tmp8983) | (tmp8982 & tmp8983);
  wire tmp8985;
  assign tmp8985 = (tmp8976 & tmp8980) | (tmp8976 & tmp8984) | (tmp8980 & tmp8984);
  wire tmp8986;
  assign tmp8986 = (tmp8959 & tmp8972) | (tmp8959 & tmp8985) | (tmp8972 & tmp8985);
  wire tmp8987;
  assign tmp8987 = (tmp8906 & tmp8946) | (tmp8906 & tmp8986) | (tmp8946 & tmp8986);
  wire tmp8988;
  assign tmp8988 = 1'b0;
  wire tmp8989;
  assign tmp8989 = 1'b0;
  wire tmp8990;
  assign tmp8990 = 1'b0;
  wire tmp8991;
  assign tmp8991 = (tmp8988 & tmp8989) | (tmp8988 & tmp8990) | (tmp8989 & tmp8990);
  wire tmp8992;
  assign tmp8992 = 1'b0;
  wire tmp8993;
  assign tmp8993 = 1'b0;
  wire tmp8994;
  assign tmp8994 = 1'b0;
  wire tmp8995;
  assign tmp8995 = (tmp8992 & tmp8993) | (tmp8992 & tmp8994) | (tmp8993 & tmp8994);
  wire tmp8996;
  assign tmp8996 = 1'b0;
  wire tmp8997;
  assign tmp8997 = 1'b0;
  wire tmp8998;
  assign tmp8998 = 1'b0;
  wire tmp8999;
  assign tmp8999 = (tmp8996 & tmp8997) | (tmp8996 & tmp8998) | (tmp8997 & tmp8998);
  wire tmp9000;
  assign tmp9000 = (tmp8991 & tmp8995) | (tmp8991 & tmp8999) | (tmp8995 & tmp8999);
  wire tmp9001;
  assign tmp9001 = 1'b0;
  wire tmp9002;
  assign tmp9002 = 1'b0;
  wire tmp9003;
  assign tmp9003 = 1'b0;
  wire tmp9004;
  assign tmp9004 = (tmp9001 & tmp9002) | (tmp9001 & tmp9003) | (tmp9002 & tmp9003);
  wire tmp9005;
  assign tmp9005 = 1'b0;
  wire tmp9006;
  assign tmp9006 = 1'b0;
  wire tmp9007;
  assign tmp9007 = 1'b0;
  wire tmp9008;
  assign tmp9008 = (tmp9005 & tmp9006) | (tmp9005 & tmp9007) | (tmp9006 & tmp9007);
  wire tmp9009;
  assign tmp9009 = 1'b0;
  wire tmp9010;
  assign tmp9010 = 1'b0;
  wire tmp9011;
  assign tmp9011 = 1'b0;
  wire tmp9012;
  assign tmp9012 = (tmp9009 & tmp9010) | (tmp9009 & tmp9011) | (tmp9010 & tmp9011);
  wire tmp9013;
  assign tmp9013 = (tmp9004 & tmp9008) | (tmp9004 & tmp9012) | (tmp9008 & tmp9012);
  wire tmp9014;
  assign tmp9014 = 1'b0;
  wire tmp9015;
  assign tmp9015 = 1'b0;
  wire tmp9016;
  assign tmp9016 = 1'b0;
  wire tmp9017;
  assign tmp9017 = (tmp9014 & tmp9015) | (tmp9014 & tmp9016) | (tmp9015 & tmp9016);
  wire tmp9018;
  assign tmp9018 = 1'b0;
  wire tmp9019;
  assign tmp9019 = 1'b0;
  wire tmp9020;
  assign tmp9020 = 1'b0;
  wire tmp9021;
  assign tmp9021 = (tmp9018 & tmp9019) | (tmp9018 & tmp9020) | (tmp9019 & tmp9020);
  wire tmp9022;
  assign tmp9022 = 1'b0;
  wire tmp9023;
  assign tmp9023 = 1'b0;
  wire tmp9024;
  assign tmp9024 = 1'b0;
  wire tmp9025;
  assign tmp9025 = (tmp9022 & tmp9023) | (tmp9022 & tmp9024) | (tmp9023 & tmp9024);
  wire tmp9026;
  assign tmp9026 = (tmp9017 & tmp9021) | (tmp9017 & tmp9025) | (tmp9021 & tmp9025);
  wire tmp9027;
  assign tmp9027 = (tmp9000 & tmp9013) | (tmp9000 & tmp9026) | (tmp9013 & tmp9026);
  wire tmp9028;
  assign tmp9028 = 1'b0;
  wire tmp9029;
  assign tmp9029 = 1'b0;
  wire tmp9030;
  assign tmp9030 = 1'b0;
  wire tmp9031;
  assign tmp9031 = (tmp9028 & tmp9029) | (tmp9028 & tmp9030) | (tmp9029 & tmp9030);
  wire tmp9032;
  assign tmp9032 = 1'b0;
  wire tmp9033;
  assign tmp9033 = 1'b0;
  wire tmp9034;
  assign tmp9034 = 1'b0;
  wire tmp9035;
  assign tmp9035 = (tmp9032 & tmp9033) | (tmp9032 & tmp9034) | (tmp9033 & tmp9034);
  wire tmp9036;
  assign tmp9036 = 1'b0;
  wire tmp9037;
  assign tmp9037 = 1'b0;
  wire tmp9038;
  assign tmp9038 = 1'b0;
  wire tmp9039;
  assign tmp9039 = (tmp9036 & tmp9037) | (tmp9036 & tmp9038) | (tmp9037 & tmp9038);
  wire tmp9040;
  assign tmp9040 = (tmp9031 & tmp9035) | (tmp9031 & tmp9039) | (tmp9035 & tmp9039);
  wire tmp9041;
  assign tmp9041 = 1'b0;
  wire tmp9042;
  assign tmp9042 = 1'b0;
  wire tmp9043;
  assign tmp9043 = 1'b0;
  wire tmp9044;
  assign tmp9044 = (tmp9041 & tmp9042) | (tmp9041 & tmp9043) | (tmp9042 & tmp9043);
  wire tmp9045;
  assign tmp9045 = 1'b0;
  wire tmp9046;
  assign tmp9046 = ~pi7;
  wire tmp9047;
  assign tmp9047 = 1'b0;
  wire tmp9048;
  assign tmp9048 = (tmp9045 & tmp9046) | (tmp9045 & tmp9047) | (tmp9046 & tmp9047);
  wire tmp9049;
  assign tmp9049 = 1'b0;
  wire tmp9050;
  assign tmp9050 = 1'b0;
  wire tmp9051;
  assign tmp9051 = 1'b0;
  wire tmp9052;
  assign tmp9052 = (tmp9049 & tmp9050) | (tmp9049 & tmp9051) | (tmp9050 & tmp9051);
  wire tmp9053;
  assign tmp9053 = (tmp9044 & tmp9048) | (tmp9044 & tmp9052) | (tmp9048 & tmp9052);
  wire tmp9054;
  assign tmp9054 = 1'b0;
  wire tmp9055;
  assign tmp9055 = 1'b0;
  wire tmp9056;
  assign tmp9056 = 1'b0;
  wire tmp9057;
  assign tmp9057 = (tmp9054 & tmp9055) | (tmp9054 & tmp9056) | (tmp9055 & tmp9056);
  wire tmp9058;
  assign tmp9058 = 1'b0;
  wire tmp9059;
  assign tmp9059 = 1'b0;
  wire tmp9060;
  assign tmp9060 = 1'b0;
  wire tmp9061;
  assign tmp9061 = (tmp9058 & tmp9059) | (tmp9058 & tmp9060) | (tmp9059 & tmp9060);
  wire tmp9062;
  assign tmp9062 = 1'b0;
  wire tmp9063;
  assign tmp9063 = 1'b0;
  wire tmp9064;
  assign tmp9064 = 1'b0;
  wire tmp9065;
  assign tmp9065 = (tmp9062 & tmp9063) | (tmp9062 & tmp9064) | (tmp9063 & tmp9064);
  wire tmp9066;
  assign tmp9066 = (tmp9057 & tmp9061) | (tmp9057 & tmp9065) | (tmp9061 & tmp9065);
  wire tmp9067;
  assign tmp9067 = (tmp9040 & tmp9053) | (tmp9040 & tmp9066) | (tmp9053 & tmp9066);
  wire tmp9068;
  assign tmp9068 = 1'b0;
  wire tmp9069;
  assign tmp9069 = 1'b0;
  wire tmp9070;
  assign tmp9070 = 1'b0;
  wire tmp9071;
  assign tmp9071 = (tmp9068 & tmp9069) | (tmp9068 & tmp9070) | (tmp9069 & tmp9070);
  wire tmp9072;
  assign tmp9072 = 1'b0;
  wire tmp9073;
  assign tmp9073 = 1'b0;
  wire tmp9074;
  assign tmp9074 = 1'b0;
  wire tmp9075;
  assign tmp9075 = (tmp9072 & tmp9073) | (tmp9072 & tmp9074) | (tmp9073 & tmp9074);
  wire tmp9076;
  assign tmp9076 = 1'b0;
  wire tmp9077;
  assign tmp9077 = 1'b0;
  wire tmp9078;
  assign tmp9078 = 1'b0;
  wire tmp9079;
  assign tmp9079 = (tmp9076 & tmp9077) | (tmp9076 & tmp9078) | (tmp9077 & tmp9078);
  wire tmp9080;
  assign tmp9080 = (tmp9071 & tmp9075) | (tmp9071 & tmp9079) | (tmp9075 & tmp9079);
  wire tmp9081;
  assign tmp9081 = 1'b0;
  wire tmp9082;
  assign tmp9082 = 1'b0;
  wire tmp9083;
  assign tmp9083 = 1'b0;
  wire tmp9084;
  assign tmp9084 = (tmp9081 & tmp9082) | (tmp9081 & tmp9083) | (tmp9082 & tmp9083);
  wire tmp9085;
  assign tmp9085 = 1'b0;
  wire tmp9086;
  assign tmp9086 = 1'b0;
  wire tmp9087;
  assign tmp9087 = 1'b0;
  wire tmp9088;
  assign tmp9088 = (tmp9085 & tmp9086) | (tmp9085 & tmp9087) | (tmp9086 & tmp9087);
  wire tmp9089;
  assign tmp9089 = 1'b0;
  wire tmp9090;
  assign tmp9090 = 1'b0;
  wire tmp9091;
  assign tmp9091 = 1'b0;
  wire tmp9092;
  assign tmp9092 = (tmp9089 & tmp9090) | (tmp9089 & tmp9091) | (tmp9090 & tmp9091);
  wire tmp9093;
  assign tmp9093 = (tmp9084 & tmp9088) | (tmp9084 & tmp9092) | (tmp9088 & tmp9092);
  wire tmp9094;
  assign tmp9094 = 1'b0;
  wire tmp9095;
  assign tmp9095 = 1'b0;
  wire tmp9096;
  assign tmp9096 = 1'b0;
  wire tmp9097;
  assign tmp9097 = (tmp9094 & tmp9095) | (tmp9094 & tmp9096) | (tmp9095 & tmp9096);
  wire tmp9098;
  assign tmp9098 = 1'b0;
  wire tmp9099;
  assign tmp9099 = 1'b0;
  wire tmp9100;
  assign tmp9100 = 1'b0;
  wire tmp9101;
  assign tmp9101 = (tmp9098 & tmp9099) | (tmp9098 & tmp9100) | (tmp9099 & tmp9100);
  wire tmp9102;
  assign tmp9102 = 1'b0;
  wire tmp9103;
  assign tmp9103 = 1'b0;
  wire tmp9104;
  assign tmp9104 = 1'b0;
  wire tmp9105;
  assign tmp9105 = (tmp9102 & tmp9103) | (tmp9102 & tmp9104) | (tmp9103 & tmp9104);
  wire tmp9106;
  assign tmp9106 = (tmp9097 & tmp9101) | (tmp9097 & tmp9105) | (tmp9101 & tmp9105);
  wire tmp9107;
  assign tmp9107 = (tmp9080 & tmp9093) | (tmp9080 & tmp9106) | (tmp9093 & tmp9106);
  wire tmp9108;
  assign tmp9108 = (tmp9027 & tmp9067) | (tmp9027 & tmp9107) | (tmp9067 & tmp9107);
  wire tmp9109;
  assign tmp9109 = (tmp8866 & tmp8987) | (tmp8866 & tmp9108) | (tmp8987 & tmp9108);
  wire tmp9110;
  assign tmp9110 = 1'b0;
  wire tmp9111;
  assign tmp9111 = 1'b0;
  wire tmp9112;
  assign tmp9112 = 1'b0;
  wire tmp9113;
  assign tmp9113 = (tmp9110 & tmp9111) | (tmp9110 & tmp9112) | (tmp9111 & tmp9112);
  wire tmp9114;
  assign tmp9114 = 1'b0;
  wire tmp9115;
  assign tmp9115 = 1'b0;
  wire tmp9116;
  assign tmp9116 = 1'b0;
  wire tmp9117;
  assign tmp9117 = (tmp9114 & tmp9115) | (tmp9114 & tmp9116) | (tmp9115 & tmp9116);
  wire tmp9118;
  assign tmp9118 = 1'b0;
  wire tmp9119;
  assign tmp9119 = 1'b0;
  wire tmp9120;
  assign tmp9120 = 1'b0;
  wire tmp9121;
  assign tmp9121 = (tmp9118 & tmp9119) | (tmp9118 & tmp9120) | (tmp9119 & tmp9120);
  wire tmp9122;
  assign tmp9122 = (tmp9113 & tmp9117) | (tmp9113 & tmp9121) | (tmp9117 & tmp9121);
  wire tmp9123;
  assign tmp9123 = 1'b0;
  wire tmp9124;
  assign tmp9124 = 1'b0;
  wire tmp9125;
  assign tmp9125 = 1'b0;
  wire tmp9126;
  assign tmp9126 = (tmp9123 & tmp9124) | (tmp9123 & tmp9125) | (tmp9124 & tmp9125);
  wire tmp9127;
  assign tmp9127 = 1'b0;
  wire tmp9128;
  assign tmp9128 = 1'b1;
  wire tmp9129;
  assign tmp9129 = 1'b0;
  wire tmp9130;
  assign tmp9130 = (tmp9127 & tmp9128) | (tmp9127 & tmp9129) | (tmp9128 & tmp9129);
  wire tmp9131;
  assign tmp9131 = 1'b0;
  wire tmp9132;
  assign tmp9132 = 1'b0;
  wire tmp9133;
  assign tmp9133 = 1'b0;
  wire tmp9134;
  assign tmp9134 = (tmp9131 & tmp9132) | (tmp9131 & tmp9133) | (tmp9132 & tmp9133);
  wire tmp9135;
  assign tmp9135 = (tmp9126 & tmp9130) | (tmp9126 & tmp9134) | (tmp9130 & tmp9134);
  wire tmp9136;
  assign tmp9136 = 1'b0;
  wire tmp9137;
  assign tmp9137 = 1'b0;
  wire tmp9138;
  assign tmp9138 = 1'b0;
  wire tmp9139;
  assign tmp9139 = (tmp9136 & tmp9137) | (tmp9136 & tmp9138) | (tmp9137 & tmp9138);
  wire tmp9140;
  assign tmp9140 = 1'b0;
  wire tmp9141;
  assign tmp9141 = 1'b0;
  wire tmp9142;
  assign tmp9142 = 1'b0;
  wire tmp9143;
  assign tmp9143 = (tmp9140 & tmp9141) | (tmp9140 & tmp9142) | (tmp9141 & tmp9142);
  wire tmp9144;
  assign tmp9144 = 1'b0;
  wire tmp9145;
  assign tmp9145 = 1'b0;
  wire tmp9146;
  assign tmp9146 = 1'b0;
  wire tmp9147;
  assign tmp9147 = (tmp9144 & tmp9145) | (tmp9144 & tmp9146) | (tmp9145 & tmp9146);
  wire tmp9148;
  assign tmp9148 = (tmp9139 & tmp9143) | (tmp9139 & tmp9147) | (tmp9143 & tmp9147);
  wire tmp9149;
  assign tmp9149 = (tmp9122 & tmp9135) | (tmp9122 & tmp9148) | (tmp9135 & tmp9148);
  wire tmp9150;
  assign tmp9150 = 1'b0;
  wire tmp9151;
  assign tmp9151 = 1'b0;
  wire tmp9152;
  assign tmp9152 = 1'b0;
  wire tmp9153;
  assign tmp9153 = (tmp9150 & tmp9151) | (tmp9150 & tmp9152) | (tmp9151 & tmp9152);
  wire tmp9154;
  assign tmp9154 = 1'b0;
  wire tmp9155;
  assign tmp9155 = 1'b1;
  wire tmp9156;
  assign tmp9156 = 1'b0;
  wire tmp9157;
  assign tmp9157 = (tmp9154 & tmp9155) | (tmp9154 & tmp9156) | (tmp9155 & tmp9156);
  wire tmp9158;
  assign tmp9158 = 1'b0;
  wire tmp9159;
  assign tmp9159 = 1'b0;
  wire tmp9160;
  assign tmp9160 = 1'b0;
  wire tmp9161;
  assign tmp9161 = (tmp9158 & tmp9159) | (tmp9158 & tmp9160) | (tmp9159 & tmp9160);
  wire tmp9162;
  assign tmp9162 = (tmp9153 & tmp9157) | (tmp9153 & tmp9161) | (tmp9157 & tmp9161);
  wire tmp9163;
  assign tmp9163 = 1'b0;
  wire tmp9164;
  assign tmp9164 = 1'b1;
  wire tmp9165;
  assign tmp9165 = 1'b0;
  wire tmp9166;
  assign tmp9166 = (tmp9163 & tmp9164) | (tmp9163 & tmp9165) | (tmp9164 & tmp9165);
  wire tmp9167;
  assign tmp9167 = 1'b1;
  wire tmp9168;
  assign tmp9168 = ~pi6;
  wire tmp9169;
  assign tmp9169 = ~pi7;
  wire tmp9170;
  assign tmp9170 = (tmp9167 & tmp9168) | (tmp9167 & tmp9169) | (tmp9168 & tmp9169);
  wire tmp9171;
  assign tmp9171 = 1'b0;
  wire tmp9172;
  assign tmp9172 = ~pi7;
  wire tmp9173;
  assign tmp9173 = 1'b0;
  wire tmp9174;
  assign tmp9174 = (tmp9171 & tmp9172) | (tmp9171 & tmp9173) | (tmp9172 & tmp9173);
  wire tmp9175;
  assign tmp9175 = (tmp9166 & tmp9170) | (tmp9166 & tmp9174) | (tmp9170 & tmp9174);
  wire tmp9176;
  assign tmp9176 = 1'b0;
  wire tmp9177;
  assign tmp9177 = 1'b0;
  wire tmp9178;
  assign tmp9178 = 1'b0;
  wire tmp9179;
  assign tmp9179 = (tmp9176 & tmp9177) | (tmp9176 & tmp9178) | (tmp9177 & tmp9178);
  wire tmp9180;
  assign tmp9180 = 1'b0;
  wire tmp9181;
  assign tmp9181 = ~pi7;
  wire tmp9182;
  assign tmp9182 = 1'b0;
  wire tmp9183;
  assign tmp9183 = (tmp9180 & tmp9181) | (tmp9180 & tmp9182) | (tmp9181 & tmp9182);
  wire tmp9184;
  assign tmp9184 = 1'b0;
  wire tmp9185;
  assign tmp9185 = 1'b0;
  wire tmp9186;
  assign tmp9186 = 1'b0;
  wire tmp9187;
  assign tmp9187 = (tmp9184 & tmp9185) | (tmp9184 & tmp9186) | (tmp9185 & tmp9186);
  wire tmp9188;
  assign tmp9188 = (tmp9179 & tmp9183) | (tmp9179 & tmp9187) | (tmp9183 & tmp9187);
  wire tmp9189;
  assign tmp9189 = (tmp9162 & tmp9175) | (tmp9162 & tmp9188) | (tmp9175 & tmp9188);
  wire tmp9190;
  assign tmp9190 = 1'b0;
  wire tmp9191;
  assign tmp9191 = 1'b0;
  wire tmp9192;
  assign tmp9192 = 1'b0;
  wire tmp9193;
  assign tmp9193 = (tmp9190 & tmp9191) | (tmp9190 & tmp9192) | (tmp9191 & tmp9192);
  wire tmp9194;
  assign tmp9194 = 1'b0;
  wire tmp9195;
  assign tmp9195 = 1'b0;
  wire tmp9196;
  assign tmp9196 = 1'b0;
  wire tmp9197;
  assign tmp9197 = (tmp9194 & tmp9195) | (tmp9194 & tmp9196) | (tmp9195 & tmp9196);
  wire tmp9198;
  assign tmp9198 = 1'b0;
  wire tmp9199;
  assign tmp9199 = 1'b0;
  wire tmp9200;
  assign tmp9200 = 1'b0;
  wire tmp9201;
  assign tmp9201 = (tmp9198 & tmp9199) | (tmp9198 & tmp9200) | (tmp9199 & tmp9200);
  wire tmp9202;
  assign tmp9202 = (tmp9193 & tmp9197) | (tmp9193 & tmp9201) | (tmp9197 & tmp9201);
  wire tmp9203;
  assign tmp9203 = 1'b0;
  wire tmp9204;
  assign tmp9204 = 1'b0;
  wire tmp9205;
  assign tmp9205 = 1'b0;
  wire tmp9206;
  assign tmp9206 = (tmp9203 & tmp9204) | (tmp9203 & tmp9205) | (tmp9204 & tmp9205);
  wire tmp9207;
  assign tmp9207 = 1'b0;
  wire tmp9208;
  assign tmp9208 = ~pi7;
  wire tmp9209;
  assign tmp9209 = 1'b0;
  wire tmp9210;
  assign tmp9210 = (tmp9207 & tmp9208) | (tmp9207 & tmp9209) | (tmp9208 & tmp9209);
  wire tmp9211;
  assign tmp9211 = 1'b0;
  wire tmp9212;
  assign tmp9212 = 1'b0;
  wire tmp9213;
  assign tmp9213 = 1'b0;
  wire tmp9214;
  assign tmp9214 = (tmp9211 & tmp9212) | (tmp9211 & tmp9213) | (tmp9212 & tmp9213);
  wire tmp9215;
  assign tmp9215 = (tmp9206 & tmp9210) | (tmp9206 & tmp9214) | (tmp9210 & tmp9214);
  wire tmp9216;
  assign tmp9216 = 1'b0;
  wire tmp9217;
  assign tmp9217 = 1'b0;
  wire tmp9218;
  assign tmp9218 = 1'b0;
  wire tmp9219;
  assign tmp9219 = (tmp9216 & tmp9217) | (tmp9216 & tmp9218) | (tmp9217 & tmp9218);
  wire tmp9220;
  assign tmp9220 = 1'b0;
  wire tmp9221;
  assign tmp9221 = 1'b0;
  wire tmp9222;
  assign tmp9222 = 1'b0;
  wire tmp9223;
  assign tmp9223 = (tmp9220 & tmp9221) | (tmp9220 & tmp9222) | (tmp9221 & tmp9222);
  wire tmp9224;
  assign tmp9224 = 1'b0;
  wire tmp9225;
  assign tmp9225 = 1'b0;
  wire tmp9226;
  assign tmp9226 = 1'b0;
  wire tmp9227;
  assign tmp9227 = (tmp9224 & tmp9225) | (tmp9224 & tmp9226) | (tmp9225 & tmp9226);
  wire tmp9228;
  assign tmp9228 = (tmp9219 & tmp9223) | (tmp9219 & tmp9227) | (tmp9223 & tmp9227);
  wire tmp9229;
  assign tmp9229 = (tmp9202 & tmp9215) | (tmp9202 & tmp9228) | (tmp9215 & tmp9228);
  wire tmp9230;
  assign tmp9230 = (tmp9149 & tmp9189) | (tmp9149 & tmp9229) | (tmp9189 & tmp9229);
  wire tmp9231;
  assign tmp9231 = 1'b0;
  wire tmp9232;
  assign tmp9232 = 1'b0;
  wire tmp9233;
  assign tmp9233 = 1'b0;
  wire tmp9234;
  assign tmp9234 = (tmp9231 & tmp9232) | (tmp9231 & tmp9233) | (tmp9232 & tmp9233);
  wire tmp9235;
  assign tmp9235 = 1'b0;
  wire tmp9236;
  assign tmp9236 = 1'b1;
  wire tmp9237;
  assign tmp9237 = 1'b0;
  wire tmp9238;
  assign tmp9238 = (tmp9235 & tmp9236) | (tmp9235 & tmp9237) | (tmp9236 & tmp9237);
  wire tmp9239;
  assign tmp9239 = 1'b0;
  wire tmp9240;
  assign tmp9240 = 1'b0;
  wire tmp9241;
  assign tmp9241 = 1'b0;
  wire tmp9242;
  assign tmp9242 = (tmp9239 & tmp9240) | (tmp9239 & tmp9241) | (tmp9240 & tmp9241);
  wire tmp9243;
  assign tmp9243 = (tmp9234 & tmp9238) | (tmp9234 & tmp9242) | (tmp9238 & tmp9242);
  wire tmp9244;
  assign tmp9244 = 1'b0;
  wire tmp9245;
  assign tmp9245 = 1'b1;
  wire tmp9246;
  assign tmp9246 = 1'b0;
  wire tmp9247;
  assign tmp9247 = (tmp9244 & tmp9245) | (tmp9244 & tmp9246) | (tmp9245 & tmp9246);
  wire tmp9248;
  assign tmp9248 = 1'b1;
  wire tmp9249;
  assign tmp9249 = ~pi6;
  wire tmp9250;
  assign tmp9250 = ~pi7;
  wire tmp9251;
  assign tmp9251 = (tmp9248 & tmp9249) | (tmp9248 & tmp9250) | (tmp9249 & tmp9250);
  wire tmp9252;
  assign tmp9252 = 1'b0;
  wire tmp9253;
  assign tmp9253 = ~pi7;
  wire tmp9254;
  assign tmp9254 = 1'b0;
  wire tmp9255;
  assign tmp9255 = (tmp9252 & tmp9253) | (tmp9252 & tmp9254) | (tmp9253 & tmp9254);
  wire tmp9256;
  assign tmp9256 = (tmp9247 & tmp9251) | (tmp9247 & tmp9255) | (tmp9251 & tmp9255);
  wire tmp9257;
  assign tmp9257 = 1'b0;
  wire tmp9258;
  assign tmp9258 = 1'b0;
  wire tmp9259;
  assign tmp9259 = 1'b0;
  wire tmp9260;
  assign tmp9260 = (tmp9257 & tmp9258) | (tmp9257 & tmp9259) | (tmp9258 & tmp9259);
  wire tmp9261;
  assign tmp9261 = 1'b0;
  wire tmp9262;
  assign tmp9262 = ~pi7;
  wire tmp9263;
  assign tmp9263 = 1'b0;
  wire tmp9264;
  assign tmp9264 = (tmp9261 & tmp9262) | (tmp9261 & tmp9263) | (tmp9262 & tmp9263);
  wire tmp9265;
  assign tmp9265 = 1'b0;
  wire tmp9266;
  assign tmp9266 = 1'b0;
  wire tmp9267;
  assign tmp9267 = 1'b0;
  wire tmp9268;
  assign tmp9268 = (tmp9265 & tmp9266) | (tmp9265 & tmp9267) | (tmp9266 & tmp9267);
  wire tmp9269;
  assign tmp9269 = (tmp9260 & tmp9264) | (tmp9260 & tmp9268) | (tmp9264 & tmp9268);
  wire tmp9270;
  assign tmp9270 = (tmp9243 & tmp9256) | (tmp9243 & tmp9269) | (tmp9256 & tmp9269);
  wire tmp9271;
  assign tmp9271 = 1'b0;
  wire tmp9272;
  assign tmp9272 = 1'b1;
  wire tmp9273;
  assign tmp9273 = 1'b0;
  wire tmp9274;
  assign tmp9274 = (tmp9271 & tmp9272) | (tmp9271 & tmp9273) | (tmp9272 & tmp9273);
  wire tmp9275;
  assign tmp9275 = 1'b1;
  wire tmp9276;
  assign tmp9276 = ~pi6;
  wire tmp9277;
  assign tmp9277 = ~pi7;
  wire tmp9278;
  assign tmp9278 = (tmp9275 & tmp9276) | (tmp9275 & tmp9277) | (tmp9276 & tmp9277);
  wire tmp9279;
  assign tmp9279 = 1'b0;
  wire tmp9280;
  assign tmp9280 = ~pi7;
  wire tmp9281;
  assign tmp9281 = 1'b0;
  wire tmp9282;
  assign tmp9282 = (tmp9279 & tmp9280) | (tmp9279 & tmp9281) | (tmp9280 & tmp9281);
  wire tmp9283;
  assign tmp9283 = (tmp9274 & tmp9278) | (tmp9274 & tmp9282) | (tmp9278 & tmp9282);
  wire tmp9284;
  assign tmp9284 = 1'b1;
  wire tmp9285;
  assign tmp9285 = ~pi6;
  wire tmp9286;
  assign tmp9286 = ~pi7;
  wire tmp9287;
  assign tmp9287 = (tmp9284 & tmp9285) | (tmp9284 & tmp9286) | (tmp9285 & tmp9286);
  wire tmp9288;
  assign tmp9288 = ~pi6;
  wire tmp9289;
  assign tmp9289 = 1'b1;
  wire tmp9290;
  assign tmp9290 = 1'b1;
  wire tmp9291;
  assign tmp9291 = (tmp9288 & tmp9289) | (tmp9288 & tmp9290) | (tmp9289 & tmp9290);
  wire tmp9292;
  assign tmp9292 = ~pi7;
  wire tmp9293;
  assign tmp9293 = 1'b1;
  wire tmp9294;
  assign tmp9294 = 1'b0;
  wire tmp9295;
  assign tmp9295 = (tmp9292 & tmp9293) | (tmp9292 & tmp9294) | (tmp9293 & tmp9294);
  wire tmp9296;
  assign tmp9296 = (tmp9287 & tmp9291) | (tmp9287 & tmp9295) | (tmp9291 & tmp9295);
  wire tmp9297;
  assign tmp9297 = 1'b0;
  wire tmp9298;
  assign tmp9298 = ~pi7;
  wire tmp9299;
  assign tmp9299 = 1'b0;
  wire tmp9300;
  assign tmp9300 = (tmp9297 & tmp9298) | (tmp9297 & tmp9299) | (tmp9298 & tmp9299);
  wire tmp9301;
  assign tmp9301 = ~pi7;
  wire tmp9302;
  assign tmp9302 = 1'b1;
  wire tmp9303;
  assign tmp9303 = 1'b0;
  wire tmp9304;
  assign tmp9304 = (tmp9301 & tmp9302) | (tmp9301 & tmp9303) | (tmp9302 & tmp9303);
  wire tmp9305;
  assign tmp9305 = 1'b0;
  wire tmp9306;
  assign tmp9306 = 1'b0;
  wire tmp9307;
  assign tmp9307 = 1'b0;
  wire tmp9308;
  assign tmp9308 = (tmp9305 & tmp9306) | (tmp9305 & tmp9307) | (tmp9306 & tmp9307);
  wire tmp9309;
  assign tmp9309 = (tmp9300 & tmp9304) | (tmp9300 & tmp9308) | (tmp9304 & tmp9308);
  wire tmp9310;
  assign tmp9310 = (tmp9283 & tmp9296) | (tmp9283 & tmp9309) | (tmp9296 & tmp9309);
  wire tmp9311;
  assign tmp9311 = 1'b0;
  wire tmp9312;
  assign tmp9312 = 1'b0;
  wire tmp9313;
  assign tmp9313 = 1'b0;
  wire tmp9314;
  assign tmp9314 = (tmp9311 & tmp9312) | (tmp9311 & tmp9313) | (tmp9312 & tmp9313);
  wire tmp9315;
  assign tmp9315 = 1'b0;
  wire tmp9316;
  assign tmp9316 = ~pi7;
  wire tmp9317;
  assign tmp9317 = 1'b0;
  wire tmp9318;
  assign tmp9318 = (tmp9315 & tmp9316) | (tmp9315 & tmp9317) | (tmp9316 & tmp9317);
  wire tmp9319;
  assign tmp9319 = 1'b0;
  wire tmp9320;
  assign tmp9320 = 1'b0;
  wire tmp9321;
  assign tmp9321 = 1'b0;
  wire tmp9322;
  assign tmp9322 = (tmp9319 & tmp9320) | (tmp9319 & tmp9321) | (tmp9320 & tmp9321);
  wire tmp9323;
  assign tmp9323 = (tmp9314 & tmp9318) | (tmp9314 & tmp9322) | (tmp9318 & tmp9322);
  wire tmp9324;
  assign tmp9324 = 1'b0;
  wire tmp9325;
  assign tmp9325 = ~pi7;
  wire tmp9326;
  assign tmp9326 = 1'b0;
  wire tmp9327;
  assign tmp9327 = (tmp9324 & tmp9325) | (tmp9324 & tmp9326) | (tmp9325 & tmp9326);
  wire tmp9328;
  assign tmp9328 = ~pi7;
  wire tmp9329;
  assign tmp9329 = 1'b1;
  wire tmp9330;
  assign tmp9330 = 1'b0;
  wire tmp9331;
  assign tmp9331 = (tmp9328 & tmp9329) | (tmp9328 & tmp9330) | (tmp9329 & tmp9330);
  wire tmp9332;
  assign tmp9332 = 1'b0;
  wire tmp9333;
  assign tmp9333 = 1'b0;
  wire tmp9334;
  assign tmp9334 = 1'b0;
  wire tmp9335;
  assign tmp9335 = (tmp9332 & tmp9333) | (tmp9332 & tmp9334) | (tmp9333 & tmp9334);
  wire tmp9336;
  assign tmp9336 = (tmp9327 & tmp9331) | (tmp9327 & tmp9335) | (tmp9331 & tmp9335);
  wire tmp9337;
  assign tmp9337 = 1'b0;
  wire tmp9338;
  assign tmp9338 = 1'b0;
  wire tmp9339;
  assign tmp9339 = 1'b0;
  wire tmp9340;
  assign tmp9340 = (tmp9337 & tmp9338) | (tmp9337 & tmp9339) | (tmp9338 & tmp9339);
  wire tmp9341;
  assign tmp9341 = 1'b0;
  wire tmp9342;
  assign tmp9342 = 1'b0;
  wire tmp9343;
  assign tmp9343 = 1'b0;
  wire tmp9344;
  assign tmp9344 = (tmp9341 & tmp9342) | (tmp9341 & tmp9343) | (tmp9342 & tmp9343);
  wire tmp9345;
  assign tmp9345 = 1'b0;
  wire tmp9346;
  assign tmp9346 = 1'b0;
  wire tmp9347;
  assign tmp9347 = 1'b0;
  wire tmp9348;
  assign tmp9348 = (tmp9345 & tmp9346) | (tmp9345 & tmp9347) | (tmp9346 & tmp9347);
  wire tmp9349;
  assign tmp9349 = (tmp9340 & tmp9344) | (tmp9340 & tmp9348) | (tmp9344 & tmp9348);
  wire tmp9350;
  assign tmp9350 = (tmp9323 & tmp9336) | (tmp9323 & tmp9349) | (tmp9336 & tmp9349);
  wire tmp9351;
  assign tmp9351 = (tmp9270 & tmp9310) | (tmp9270 & tmp9350) | (tmp9310 & tmp9350);
  wire tmp9352;
  assign tmp9352 = 1'b0;
  wire tmp9353;
  assign tmp9353 = 1'b0;
  wire tmp9354;
  assign tmp9354 = 1'b0;
  wire tmp9355;
  assign tmp9355 = (tmp9352 & tmp9353) | (tmp9352 & tmp9354) | (tmp9353 & tmp9354);
  wire tmp9356;
  assign tmp9356 = 1'b0;
  wire tmp9357;
  assign tmp9357 = 1'b0;
  wire tmp9358;
  assign tmp9358 = 1'b0;
  wire tmp9359;
  assign tmp9359 = (tmp9356 & tmp9357) | (tmp9356 & tmp9358) | (tmp9357 & tmp9358);
  wire tmp9360;
  assign tmp9360 = 1'b0;
  wire tmp9361;
  assign tmp9361 = 1'b0;
  wire tmp9362;
  assign tmp9362 = 1'b0;
  wire tmp9363;
  assign tmp9363 = (tmp9360 & tmp9361) | (tmp9360 & tmp9362) | (tmp9361 & tmp9362);
  wire tmp9364;
  assign tmp9364 = (tmp9355 & tmp9359) | (tmp9355 & tmp9363) | (tmp9359 & tmp9363);
  wire tmp9365;
  assign tmp9365 = 1'b0;
  wire tmp9366;
  assign tmp9366 = 1'b0;
  wire tmp9367;
  assign tmp9367 = 1'b0;
  wire tmp9368;
  assign tmp9368 = (tmp9365 & tmp9366) | (tmp9365 & tmp9367) | (tmp9366 & tmp9367);
  wire tmp9369;
  assign tmp9369 = 1'b0;
  wire tmp9370;
  assign tmp9370 = ~pi7;
  wire tmp9371;
  assign tmp9371 = 1'b0;
  wire tmp9372;
  assign tmp9372 = (tmp9369 & tmp9370) | (tmp9369 & tmp9371) | (tmp9370 & tmp9371);
  wire tmp9373;
  assign tmp9373 = 1'b0;
  wire tmp9374;
  assign tmp9374 = 1'b0;
  wire tmp9375;
  assign tmp9375 = 1'b0;
  wire tmp9376;
  assign tmp9376 = (tmp9373 & tmp9374) | (tmp9373 & tmp9375) | (tmp9374 & tmp9375);
  wire tmp9377;
  assign tmp9377 = (tmp9368 & tmp9372) | (tmp9368 & tmp9376) | (tmp9372 & tmp9376);
  wire tmp9378;
  assign tmp9378 = 1'b0;
  wire tmp9379;
  assign tmp9379 = 1'b0;
  wire tmp9380;
  assign tmp9380 = 1'b0;
  wire tmp9381;
  assign tmp9381 = (tmp9378 & tmp9379) | (tmp9378 & tmp9380) | (tmp9379 & tmp9380);
  wire tmp9382;
  assign tmp9382 = 1'b0;
  wire tmp9383;
  assign tmp9383 = 1'b0;
  wire tmp9384;
  assign tmp9384 = 1'b0;
  wire tmp9385;
  assign tmp9385 = (tmp9382 & tmp9383) | (tmp9382 & tmp9384) | (tmp9383 & tmp9384);
  wire tmp9386;
  assign tmp9386 = 1'b0;
  wire tmp9387;
  assign tmp9387 = 1'b0;
  wire tmp9388;
  assign tmp9388 = 1'b0;
  wire tmp9389;
  assign tmp9389 = (tmp9386 & tmp9387) | (tmp9386 & tmp9388) | (tmp9387 & tmp9388);
  wire tmp9390;
  assign tmp9390 = (tmp9381 & tmp9385) | (tmp9381 & tmp9389) | (tmp9385 & tmp9389);
  wire tmp9391;
  assign tmp9391 = (tmp9364 & tmp9377) | (tmp9364 & tmp9390) | (tmp9377 & tmp9390);
  wire tmp9392;
  assign tmp9392 = 1'b0;
  wire tmp9393;
  assign tmp9393 = 1'b0;
  wire tmp9394;
  assign tmp9394 = 1'b0;
  wire tmp9395;
  assign tmp9395 = (tmp9392 & tmp9393) | (tmp9392 & tmp9394) | (tmp9393 & tmp9394);
  wire tmp9396;
  assign tmp9396 = 1'b0;
  wire tmp9397;
  assign tmp9397 = ~pi7;
  wire tmp9398;
  assign tmp9398 = 1'b0;
  wire tmp9399;
  assign tmp9399 = (tmp9396 & tmp9397) | (tmp9396 & tmp9398) | (tmp9397 & tmp9398);
  wire tmp9400;
  assign tmp9400 = 1'b0;
  wire tmp9401;
  assign tmp9401 = 1'b0;
  wire tmp9402;
  assign tmp9402 = 1'b0;
  wire tmp9403;
  assign tmp9403 = (tmp9400 & tmp9401) | (tmp9400 & tmp9402) | (tmp9401 & tmp9402);
  wire tmp9404;
  assign tmp9404 = (tmp9395 & tmp9399) | (tmp9395 & tmp9403) | (tmp9399 & tmp9403);
  wire tmp9405;
  assign tmp9405 = 1'b0;
  wire tmp9406;
  assign tmp9406 = ~pi7;
  wire tmp9407;
  assign tmp9407 = 1'b0;
  wire tmp9408;
  assign tmp9408 = (tmp9405 & tmp9406) | (tmp9405 & tmp9407) | (tmp9406 & tmp9407);
  wire tmp9409;
  assign tmp9409 = ~pi7;
  wire tmp9410;
  assign tmp9410 = 1'b1;
  wire tmp9411;
  assign tmp9411 = 1'b0;
  wire tmp9412;
  assign tmp9412 = (tmp9409 & tmp9410) | (tmp9409 & tmp9411) | (tmp9410 & tmp9411);
  wire tmp9413;
  assign tmp9413 = 1'b0;
  wire tmp9414;
  assign tmp9414 = 1'b0;
  wire tmp9415;
  assign tmp9415 = 1'b0;
  wire tmp9416;
  assign tmp9416 = (tmp9413 & tmp9414) | (tmp9413 & tmp9415) | (tmp9414 & tmp9415);
  wire tmp9417;
  assign tmp9417 = (tmp9408 & tmp9412) | (tmp9408 & tmp9416) | (tmp9412 & tmp9416);
  wire tmp9418;
  assign tmp9418 = 1'b0;
  wire tmp9419;
  assign tmp9419 = 1'b0;
  wire tmp9420;
  assign tmp9420 = 1'b0;
  wire tmp9421;
  assign tmp9421 = (tmp9418 & tmp9419) | (tmp9418 & tmp9420) | (tmp9419 & tmp9420);
  wire tmp9422;
  assign tmp9422 = 1'b0;
  wire tmp9423;
  assign tmp9423 = 1'b0;
  wire tmp9424;
  assign tmp9424 = 1'b0;
  wire tmp9425;
  assign tmp9425 = (tmp9422 & tmp9423) | (tmp9422 & tmp9424) | (tmp9423 & tmp9424);
  wire tmp9426;
  assign tmp9426 = 1'b0;
  wire tmp9427;
  assign tmp9427 = 1'b0;
  wire tmp9428;
  assign tmp9428 = 1'b0;
  wire tmp9429;
  assign tmp9429 = (tmp9426 & tmp9427) | (tmp9426 & tmp9428) | (tmp9427 & tmp9428);
  wire tmp9430;
  assign tmp9430 = (tmp9421 & tmp9425) | (tmp9421 & tmp9429) | (tmp9425 & tmp9429);
  wire tmp9431;
  assign tmp9431 = (tmp9404 & tmp9417) | (tmp9404 & tmp9430) | (tmp9417 & tmp9430);
  wire tmp9432;
  assign tmp9432 = 1'b0;
  wire tmp9433;
  assign tmp9433 = 1'b0;
  wire tmp9434;
  assign tmp9434 = 1'b0;
  wire tmp9435;
  assign tmp9435 = (tmp9432 & tmp9433) | (tmp9432 & tmp9434) | (tmp9433 & tmp9434);
  wire tmp9436;
  assign tmp9436 = 1'b0;
  wire tmp9437;
  assign tmp9437 = 1'b0;
  wire tmp9438;
  assign tmp9438 = 1'b0;
  wire tmp9439;
  assign tmp9439 = (tmp9436 & tmp9437) | (tmp9436 & tmp9438) | (tmp9437 & tmp9438);
  wire tmp9440;
  assign tmp9440 = 1'b0;
  wire tmp9441;
  assign tmp9441 = 1'b0;
  wire tmp9442;
  assign tmp9442 = 1'b0;
  wire tmp9443;
  assign tmp9443 = (tmp9440 & tmp9441) | (tmp9440 & tmp9442) | (tmp9441 & tmp9442);
  wire tmp9444;
  assign tmp9444 = (tmp9435 & tmp9439) | (tmp9435 & tmp9443) | (tmp9439 & tmp9443);
  wire tmp9445;
  assign tmp9445 = 1'b0;
  wire tmp9446;
  assign tmp9446 = 1'b0;
  wire tmp9447;
  assign tmp9447 = 1'b0;
  wire tmp9448;
  assign tmp9448 = (tmp9445 & tmp9446) | (tmp9445 & tmp9447) | (tmp9446 & tmp9447);
  wire tmp9449;
  assign tmp9449 = 1'b0;
  wire tmp9450;
  assign tmp9450 = 1'b0;
  wire tmp9451;
  assign tmp9451 = 1'b0;
  wire tmp9452;
  assign tmp9452 = (tmp9449 & tmp9450) | (tmp9449 & tmp9451) | (tmp9450 & tmp9451);
  wire tmp9453;
  assign tmp9453 = 1'b0;
  wire tmp9454;
  assign tmp9454 = 1'b0;
  wire tmp9455;
  assign tmp9455 = 1'b0;
  wire tmp9456;
  assign tmp9456 = (tmp9453 & tmp9454) | (tmp9453 & tmp9455) | (tmp9454 & tmp9455);
  wire tmp9457;
  assign tmp9457 = (tmp9448 & tmp9452) | (tmp9448 & tmp9456) | (tmp9452 & tmp9456);
  wire tmp9458;
  assign tmp9458 = 1'b0;
  wire tmp9459;
  assign tmp9459 = 1'b0;
  wire tmp9460;
  assign tmp9460 = 1'b0;
  wire tmp9461;
  assign tmp9461 = (tmp9458 & tmp9459) | (tmp9458 & tmp9460) | (tmp9459 & tmp9460);
  wire tmp9462;
  assign tmp9462 = 1'b0;
  wire tmp9463;
  assign tmp9463 = 1'b0;
  wire tmp9464;
  assign tmp9464 = 1'b0;
  wire tmp9465;
  assign tmp9465 = (tmp9462 & tmp9463) | (tmp9462 & tmp9464) | (tmp9463 & tmp9464);
  wire tmp9466;
  assign tmp9466 = 1'b0;
  wire tmp9467;
  assign tmp9467 = 1'b0;
  wire tmp9468;
  assign tmp9468 = 1'b0;
  wire tmp9469;
  assign tmp9469 = (tmp9466 & tmp9467) | (tmp9466 & tmp9468) | (tmp9467 & tmp9468);
  wire tmp9470;
  assign tmp9470 = (tmp9461 & tmp9465) | (tmp9461 & tmp9469) | (tmp9465 & tmp9469);
  wire tmp9471;
  assign tmp9471 = (tmp9444 & tmp9457) | (tmp9444 & tmp9470) | (tmp9457 & tmp9470);
  wire tmp9472;
  assign tmp9472 = (tmp9391 & tmp9431) | (tmp9391 & tmp9471) | (tmp9431 & tmp9471);
  wire tmp9473;
  assign tmp9473 = (tmp9230 & tmp9351) | (tmp9230 & tmp9472) | (tmp9351 & tmp9472);
  wire tmp9474;
  assign tmp9474 = 1'b0;
  wire tmp9475;
  assign tmp9475 = 1'b0;
  wire tmp9476;
  assign tmp9476 = 1'b0;
  wire tmp9477;
  assign tmp9477 = (tmp9474 & tmp9475) | (tmp9474 & tmp9476) | (tmp9475 & tmp9476);
  wire tmp9478;
  assign tmp9478 = 1'b0;
  wire tmp9479;
  assign tmp9479 = 1'b0;
  wire tmp9480;
  assign tmp9480 = 1'b0;
  wire tmp9481;
  assign tmp9481 = (tmp9478 & tmp9479) | (tmp9478 & tmp9480) | (tmp9479 & tmp9480);
  wire tmp9482;
  assign tmp9482 = 1'b0;
  wire tmp9483;
  assign tmp9483 = 1'b0;
  wire tmp9484;
  assign tmp9484 = 1'b0;
  wire tmp9485;
  assign tmp9485 = (tmp9482 & tmp9483) | (tmp9482 & tmp9484) | (tmp9483 & tmp9484);
  wire tmp9486;
  assign tmp9486 = (tmp9477 & tmp9481) | (tmp9477 & tmp9485) | (tmp9481 & tmp9485);
  wire tmp9487;
  assign tmp9487 = 1'b0;
  wire tmp9488;
  assign tmp9488 = 1'b0;
  wire tmp9489;
  assign tmp9489 = 1'b0;
  wire tmp9490;
  assign tmp9490 = (tmp9487 & tmp9488) | (tmp9487 & tmp9489) | (tmp9488 & tmp9489);
  wire tmp9491;
  assign tmp9491 = 1'b0;
  wire tmp9492;
  assign tmp9492 = 1'b0;
  wire tmp9493;
  assign tmp9493 = 1'b0;
  wire tmp9494;
  assign tmp9494 = (tmp9491 & tmp9492) | (tmp9491 & tmp9493) | (tmp9492 & tmp9493);
  wire tmp9495;
  assign tmp9495 = 1'b0;
  wire tmp9496;
  assign tmp9496 = 1'b0;
  wire tmp9497;
  assign tmp9497 = 1'b0;
  wire tmp9498;
  assign tmp9498 = (tmp9495 & tmp9496) | (tmp9495 & tmp9497) | (tmp9496 & tmp9497);
  wire tmp9499;
  assign tmp9499 = (tmp9490 & tmp9494) | (tmp9490 & tmp9498) | (tmp9494 & tmp9498);
  wire tmp9500;
  assign tmp9500 = 1'b0;
  wire tmp9501;
  assign tmp9501 = 1'b0;
  wire tmp9502;
  assign tmp9502 = 1'b0;
  wire tmp9503;
  assign tmp9503 = (tmp9500 & tmp9501) | (tmp9500 & tmp9502) | (tmp9501 & tmp9502);
  wire tmp9504;
  assign tmp9504 = 1'b0;
  wire tmp9505;
  assign tmp9505 = 1'b0;
  wire tmp9506;
  assign tmp9506 = 1'b0;
  wire tmp9507;
  assign tmp9507 = (tmp9504 & tmp9505) | (tmp9504 & tmp9506) | (tmp9505 & tmp9506);
  wire tmp9508;
  assign tmp9508 = 1'b0;
  wire tmp9509;
  assign tmp9509 = 1'b0;
  wire tmp9510;
  assign tmp9510 = 1'b0;
  wire tmp9511;
  assign tmp9511 = (tmp9508 & tmp9509) | (tmp9508 & tmp9510) | (tmp9509 & tmp9510);
  wire tmp9512;
  assign tmp9512 = (tmp9503 & tmp9507) | (tmp9503 & tmp9511) | (tmp9507 & tmp9511);
  wire tmp9513;
  assign tmp9513 = (tmp9486 & tmp9499) | (tmp9486 & tmp9512) | (tmp9499 & tmp9512);
  wire tmp9514;
  assign tmp9514 = 1'b0;
  wire tmp9515;
  assign tmp9515 = 1'b0;
  wire tmp9516;
  assign tmp9516 = 1'b0;
  wire tmp9517;
  assign tmp9517 = (tmp9514 & tmp9515) | (tmp9514 & tmp9516) | (tmp9515 & tmp9516);
  wire tmp9518;
  assign tmp9518 = 1'b0;
  wire tmp9519;
  assign tmp9519 = 1'b0;
  wire tmp9520;
  assign tmp9520 = 1'b0;
  wire tmp9521;
  assign tmp9521 = (tmp9518 & tmp9519) | (tmp9518 & tmp9520) | (tmp9519 & tmp9520);
  wire tmp9522;
  assign tmp9522 = 1'b0;
  wire tmp9523;
  assign tmp9523 = 1'b0;
  wire tmp9524;
  assign tmp9524 = 1'b0;
  wire tmp9525;
  assign tmp9525 = (tmp9522 & tmp9523) | (tmp9522 & tmp9524) | (tmp9523 & tmp9524);
  wire tmp9526;
  assign tmp9526 = (tmp9517 & tmp9521) | (tmp9517 & tmp9525) | (tmp9521 & tmp9525);
  wire tmp9527;
  assign tmp9527 = 1'b0;
  wire tmp9528;
  assign tmp9528 = 1'b0;
  wire tmp9529;
  assign tmp9529 = 1'b0;
  wire tmp9530;
  assign tmp9530 = (tmp9527 & tmp9528) | (tmp9527 & tmp9529) | (tmp9528 & tmp9529);
  wire tmp9531;
  assign tmp9531 = 1'b0;
  wire tmp9532;
  assign tmp9532 = ~pi7;
  wire tmp9533;
  assign tmp9533 = 1'b0;
  wire tmp9534;
  assign tmp9534 = (tmp9531 & tmp9532) | (tmp9531 & tmp9533) | (tmp9532 & tmp9533);
  wire tmp9535;
  assign tmp9535 = 1'b0;
  wire tmp9536;
  assign tmp9536 = 1'b0;
  wire tmp9537;
  assign tmp9537 = 1'b0;
  wire tmp9538;
  assign tmp9538 = (tmp9535 & tmp9536) | (tmp9535 & tmp9537) | (tmp9536 & tmp9537);
  wire tmp9539;
  assign tmp9539 = (tmp9530 & tmp9534) | (tmp9530 & tmp9538) | (tmp9534 & tmp9538);
  wire tmp9540;
  assign tmp9540 = 1'b0;
  wire tmp9541;
  assign tmp9541 = 1'b0;
  wire tmp9542;
  assign tmp9542 = 1'b0;
  wire tmp9543;
  assign tmp9543 = (tmp9540 & tmp9541) | (tmp9540 & tmp9542) | (tmp9541 & tmp9542);
  wire tmp9544;
  assign tmp9544 = 1'b0;
  wire tmp9545;
  assign tmp9545 = 1'b0;
  wire tmp9546;
  assign tmp9546 = 1'b0;
  wire tmp9547;
  assign tmp9547 = (tmp9544 & tmp9545) | (tmp9544 & tmp9546) | (tmp9545 & tmp9546);
  wire tmp9548;
  assign tmp9548 = 1'b0;
  wire tmp9549;
  assign tmp9549 = 1'b0;
  wire tmp9550;
  assign tmp9550 = 1'b0;
  wire tmp9551;
  assign tmp9551 = (tmp9548 & tmp9549) | (tmp9548 & tmp9550) | (tmp9549 & tmp9550);
  wire tmp9552;
  assign tmp9552 = (tmp9543 & tmp9547) | (tmp9543 & tmp9551) | (tmp9547 & tmp9551);
  wire tmp9553;
  assign tmp9553 = (tmp9526 & tmp9539) | (tmp9526 & tmp9552) | (tmp9539 & tmp9552);
  wire tmp9554;
  assign tmp9554 = 1'b0;
  wire tmp9555;
  assign tmp9555 = 1'b0;
  wire tmp9556;
  assign tmp9556 = 1'b0;
  wire tmp9557;
  assign tmp9557 = (tmp9554 & tmp9555) | (tmp9554 & tmp9556) | (tmp9555 & tmp9556);
  wire tmp9558;
  assign tmp9558 = 1'b0;
  wire tmp9559;
  assign tmp9559 = 1'b0;
  wire tmp9560;
  assign tmp9560 = 1'b0;
  wire tmp9561;
  assign tmp9561 = (tmp9558 & tmp9559) | (tmp9558 & tmp9560) | (tmp9559 & tmp9560);
  wire tmp9562;
  assign tmp9562 = 1'b0;
  wire tmp9563;
  assign tmp9563 = 1'b0;
  wire tmp9564;
  assign tmp9564 = 1'b0;
  wire tmp9565;
  assign tmp9565 = (tmp9562 & tmp9563) | (tmp9562 & tmp9564) | (tmp9563 & tmp9564);
  wire tmp9566;
  assign tmp9566 = (tmp9557 & tmp9561) | (tmp9557 & tmp9565) | (tmp9561 & tmp9565);
  wire tmp9567;
  assign tmp9567 = 1'b0;
  wire tmp9568;
  assign tmp9568 = 1'b0;
  wire tmp9569;
  assign tmp9569 = 1'b0;
  wire tmp9570;
  assign tmp9570 = (tmp9567 & tmp9568) | (tmp9567 & tmp9569) | (tmp9568 & tmp9569);
  wire tmp9571;
  assign tmp9571 = 1'b0;
  wire tmp9572;
  assign tmp9572 = 1'b0;
  wire tmp9573;
  assign tmp9573 = 1'b0;
  wire tmp9574;
  assign tmp9574 = (tmp9571 & tmp9572) | (tmp9571 & tmp9573) | (tmp9572 & tmp9573);
  wire tmp9575;
  assign tmp9575 = 1'b0;
  wire tmp9576;
  assign tmp9576 = 1'b0;
  wire tmp9577;
  assign tmp9577 = 1'b0;
  wire tmp9578;
  assign tmp9578 = (tmp9575 & tmp9576) | (tmp9575 & tmp9577) | (tmp9576 & tmp9577);
  wire tmp9579;
  assign tmp9579 = (tmp9570 & tmp9574) | (tmp9570 & tmp9578) | (tmp9574 & tmp9578);
  wire tmp9580;
  assign tmp9580 = 1'b0;
  wire tmp9581;
  assign tmp9581 = 1'b0;
  wire tmp9582;
  assign tmp9582 = 1'b0;
  wire tmp9583;
  assign tmp9583 = (tmp9580 & tmp9581) | (tmp9580 & tmp9582) | (tmp9581 & tmp9582);
  wire tmp9584;
  assign tmp9584 = 1'b0;
  wire tmp9585;
  assign tmp9585 = 1'b0;
  wire tmp9586;
  assign tmp9586 = 1'b0;
  wire tmp9587;
  assign tmp9587 = (tmp9584 & tmp9585) | (tmp9584 & tmp9586) | (tmp9585 & tmp9586);
  wire tmp9588;
  assign tmp9588 = 1'b0;
  wire tmp9589;
  assign tmp9589 = 1'b0;
  wire tmp9590;
  assign tmp9590 = 1'b0;
  wire tmp9591;
  assign tmp9591 = (tmp9588 & tmp9589) | (tmp9588 & tmp9590) | (tmp9589 & tmp9590);
  wire tmp9592;
  assign tmp9592 = (tmp9583 & tmp9587) | (tmp9583 & tmp9591) | (tmp9587 & tmp9591);
  wire tmp9593;
  assign tmp9593 = (tmp9566 & tmp9579) | (tmp9566 & tmp9592) | (tmp9579 & tmp9592);
  wire tmp9594;
  assign tmp9594 = (tmp9513 & tmp9553) | (tmp9513 & tmp9593) | (tmp9553 & tmp9593);
  wire tmp9595;
  assign tmp9595 = 1'b0;
  wire tmp9596;
  assign tmp9596 = 1'b0;
  wire tmp9597;
  assign tmp9597 = 1'b0;
  wire tmp9598;
  assign tmp9598 = (tmp9595 & tmp9596) | (tmp9595 & tmp9597) | (tmp9596 & tmp9597);
  wire tmp9599;
  assign tmp9599 = 1'b0;
  wire tmp9600;
  assign tmp9600 = 1'b0;
  wire tmp9601;
  assign tmp9601 = 1'b0;
  wire tmp9602;
  assign tmp9602 = (tmp9599 & tmp9600) | (tmp9599 & tmp9601) | (tmp9600 & tmp9601);
  wire tmp9603;
  assign tmp9603 = 1'b0;
  wire tmp9604;
  assign tmp9604 = 1'b0;
  wire tmp9605;
  assign tmp9605 = 1'b0;
  wire tmp9606;
  assign tmp9606 = (tmp9603 & tmp9604) | (tmp9603 & tmp9605) | (tmp9604 & tmp9605);
  wire tmp9607;
  assign tmp9607 = (tmp9598 & tmp9602) | (tmp9598 & tmp9606) | (tmp9602 & tmp9606);
  wire tmp9608;
  assign tmp9608 = 1'b0;
  wire tmp9609;
  assign tmp9609 = 1'b0;
  wire tmp9610;
  assign tmp9610 = 1'b0;
  wire tmp9611;
  assign tmp9611 = (tmp9608 & tmp9609) | (tmp9608 & tmp9610) | (tmp9609 & tmp9610);
  wire tmp9612;
  assign tmp9612 = 1'b0;
  wire tmp9613;
  assign tmp9613 = ~pi7;
  wire tmp9614;
  assign tmp9614 = 1'b0;
  wire tmp9615;
  assign tmp9615 = (tmp9612 & tmp9613) | (tmp9612 & tmp9614) | (tmp9613 & tmp9614);
  wire tmp9616;
  assign tmp9616 = 1'b0;
  wire tmp9617;
  assign tmp9617 = 1'b0;
  wire tmp9618;
  assign tmp9618 = 1'b0;
  wire tmp9619;
  assign tmp9619 = (tmp9616 & tmp9617) | (tmp9616 & tmp9618) | (tmp9617 & tmp9618);
  wire tmp9620;
  assign tmp9620 = (tmp9611 & tmp9615) | (tmp9611 & tmp9619) | (tmp9615 & tmp9619);
  wire tmp9621;
  assign tmp9621 = 1'b0;
  wire tmp9622;
  assign tmp9622 = 1'b0;
  wire tmp9623;
  assign tmp9623 = 1'b0;
  wire tmp9624;
  assign tmp9624 = (tmp9621 & tmp9622) | (tmp9621 & tmp9623) | (tmp9622 & tmp9623);
  wire tmp9625;
  assign tmp9625 = 1'b0;
  wire tmp9626;
  assign tmp9626 = 1'b0;
  wire tmp9627;
  assign tmp9627 = 1'b0;
  wire tmp9628;
  assign tmp9628 = (tmp9625 & tmp9626) | (tmp9625 & tmp9627) | (tmp9626 & tmp9627);
  wire tmp9629;
  assign tmp9629 = 1'b0;
  wire tmp9630;
  assign tmp9630 = 1'b0;
  wire tmp9631;
  assign tmp9631 = 1'b0;
  wire tmp9632;
  assign tmp9632 = (tmp9629 & tmp9630) | (tmp9629 & tmp9631) | (tmp9630 & tmp9631);
  wire tmp9633;
  assign tmp9633 = (tmp9624 & tmp9628) | (tmp9624 & tmp9632) | (tmp9628 & tmp9632);
  wire tmp9634;
  assign tmp9634 = (tmp9607 & tmp9620) | (tmp9607 & tmp9633) | (tmp9620 & tmp9633);
  wire tmp9635;
  assign tmp9635 = 1'b0;
  wire tmp9636;
  assign tmp9636 = 1'b0;
  wire tmp9637;
  assign tmp9637 = 1'b0;
  wire tmp9638;
  assign tmp9638 = (tmp9635 & tmp9636) | (tmp9635 & tmp9637) | (tmp9636 & tmp9637);
  wire tmp9639;
  assign tmp9639 = 1'b0;
  wire tmp9640;
  assign tmp9640 = ~pi7;
  wire tmp9641;
  assign tmp9641 = 1'b0;
  wire tmp9642;
  assign tmp9642 = (tmp9639 & tmp9640) | (tmp9639 & tmp9641) | (tmp9640 & tmp9641);
  wire tmp9643;
  assign tmp9643 = 1'b0;
  wire tmp9644;
  assign tmp9644 = 1'b0;
  wire tmp9645;
  assign tmp9645 = 1'b0;
  wire tmp9646;
  assign tmp9646 = (tmp9643 & tmp9644) | (tmp9643 & tmp9645) | (tmp9644 & tmp9645);
  wire tmp9647;
  assign tmp9647 = (tmp9638 & tmp9642) | (tmp9638 & tmp9646) | (tmp9642 & tmp9646);
  wire tmp9648;
  assign tmp9648 = 1'b0;
  wire tmp9649;
  assign tmp9649 = ~pi7;
  wire tmp9650;
  assign tmp9650 = 1'b0;
  wire tmp9651;
  assign tmp9651 = (tmp9648 & tmp9649) | (tmp9648 & tmp9650) | (tmp9649 & tmp9650);
  wire tmp9652;
  assign tmp9652 = ~pi7;
  wire tmp9653;
  assign tmp9653 = 1'b1;
  wire tmp9654;
  assign tmp9654 = 1'b0;
  wire tmp9655;
  assign tmp9655 = (tmp9652 & tmp9653) | (tmp9652 & tmp9654) | (tmp9653 & tmp9654);
  wire tmp9656;
  assign tmp9656 = 1'b0;
  wire tmp9657;
  assign tmp9657 = 1'b0;
  wire tmp9658;
  assign tmp9658 = 1'b0;
  wire tmp9659;
  assign tmp9659 = (tmp9656 & tmp9657) | (tmp9656 & tmp9658) | (tmp9657 & tmp9658);
  wire tmp9660;
  assign tmp9660 = (tmp9651 & tmp9655) | (tmp9651 & tmp9659) | (tmp9655 & tmp9659);
  wire tmp9661;
  assign tmp9661 = 1'b0;
  wire tmp9662;
  assign tmp9662 = 1'b0;
  wire tmp9663;
  assign tmp9663 = 1'b0;
  wire tmp9664;
  assign tmp9664 = (tmp9661 & tmp9662) | (tmp9661 & tmp9663) | (tmp9662 & tmp9663);
  wire tmp9665;
  assign tmp9665 = 1'b0;
  wire tmp9666;
  assign tmp9666 = 1'b0;
  wire tmp9667;
  assign tmp9667 = 1'b0;
  wire tmp9668;
  assign tmp9668 = (tmp9665 & tmp9666) | (tmp9665 & tmp9667) | (tmp9666 & tmp9667);
  wire tmp9669;
  assign tmp9669 = 1'b0;
  wire tmp9670;
  assign tmp9670 = 1'b0;
  wire tmp9671;
  assign tmp9671 = 1'b0;
  wire tmp9672;
  assign tmp9672 = (tmp9669 & tmp9670) | (tmp9669 & tmp9671) | (tmp9670 & tmp9671);
  wire tmp9673;
  assign tmp9673 = (tmp9664 & tmp9668) | (tmp9664 & tmp9672) | (tmp9668 & tmp9672);
  wire tmp9674;
  assign tmp9674 = (tmp9647 & tmp9660) | (tmp9647 & tmp9673) | (tmp9660 & tmp9673);
  wire tmp9675;
  assign tmp9675 = 1'b0;
  wire tmp9676;
  assign tmp9676 = 1'b0;
  wire tmp9677;
  assign tmp9677 = 1'b0;
  wire tmp9678;
  assign tmp9678 = (tmp9675 & tmp9676) | (tmp9675 & tmp9677) | (tmp9676 & tmp9677);
  wire tmp9679;
  assign tmp9679 = 1'b0;
  wire tmp9680;
  assign tmp9680 = 1'b0;
  wire tmp9681;
  assign tmp9681 = 1'b0;
  wire tmp9682;
  assign tmp9682 = (tmp9679 & tmp9680) | (tmp9679 & tmp9681) | (tmp9680 & tmp9681);
  wire tmp9683;
  assign tmp9683 = 1'b0;
  wire tmp9684;
  assign tmp9684 = 1'b0;
  wire tmp9685;
  assign tmp9685 = 1'b0;
  wire tmp9686;
  assign tmp9686 = (tmp9683 & tmp9684) | (tmp9683 & tmp9685) | (tmp9684 & tmp9685);
  wire tmp9687;
  assign tmp9687 = (tmp9678 & tmp9682) | (tmp9678 & tmp9686) | (tmp9682 & tmp9686);
  wire tmp9688;
  assign tmp9688 = 1'b0;
  wire tmp9689;
  assign tmp9689 = 1'b0;
  wire tmp9690;
  assign tmp9690 = 1'b0;
  wire tmp9691;
  assign tmp9691 = (tmp9688 & tmp9689) | (tmp9688 & tmp9690) | (tmp9689 & tmp9690);
  wire tmp9692;
  assign tmp9692 = 1'b0;
  wire tmp9693;
  assign tmp9693 = 1'b0;
  wire tmp9694;
  assign tmp9694 = 1'b0;
  wire tmp9695;
  assign tmp9695 = (tmp9692 & tmp9693) | (tmp9692 & tmp9694) | (tmp9693 & tmp9694);
  wire tmp9696;
  assign tmp9696 = 1'b0;
  wire tmp9697;
  assign tmp9697 = 1'b0;
  wire tmp9698;
  assign tmp9698 = 1'b0;
  wire tmp9699;
  assign tmp9699 = (tmp9696 & tmp9697) | (tmp9696 & tmp9698) | (tmp9697 & tmp9698);
  wire tmp9700;
  assign tmp9700 = (tmp9691 & tmp9695) | (tmp9691 & tmp9699) | (tmp9695 & tmp9699);
  wire tmp9701;
  assign tmp9701 = 1'b0;
  wire tmp9702;
  assign tmp9702 = 1'b0;
  wire tmp9703;
  assign tmp9703 = 1'b0;
  wire tmp9704;
  assign tmp9704 = (tmp9701 & tmp9702) | (tmp9701 & tmp9703) | (tmp9702 & tmp9703);
  wire tmp9705;
  assign tmp9705 = 1'b0;
  wire tmp9706;
  assign tmp9706 = 1'b0;
  wire tmp9707;
  assign tmp9707 = 1'b0;
  wire tmp9708;
  assign tmp9708 = (tmp9705 & tmp9706) | (tmp9705 & tmp9707) | (tmp9706 & tmp9707);
  wire tmp9709;
  assign tmp9709 = 1'b0;
  wire tmp9710;
  assign tmp9710 = 1'b0;
  wire tmp9711;
  assign tmp9711 = 1'b0;
  wire tmp9712;
  assign tmp9712 = (tmp9709 & tmp9710) | (tmp9709 & tmp9711) | (tmp9710 & tmp9711);
  wire tmp9713;
  assign tmp9713 = (tmp9704 & tmp9708) | (tmp9704 & tmp9712) | (tmp9708 & tmp9712);
  wire tmp9714;
  assign tmp9714 = (tmp9687 & tmp9700) | (tmp9687 & tmp9713) | (tmp9700 & tmp9713);
  wire tmp9715;
  assign tmp9715 = (tmp9634 & tmp9674) | (tmp9634 & tmp9714) | (tmp9674 & tmp9714);
  wire tmp9716;
  assign tmp9716 = 1'b0;
  wire tmp9717;
  assign tmp9717 = 1'b0;
  wire tmp9718;
  assign tmp9718 = 1'b0;
  wire tmp9719;
  assign tmp9719 = (tmp9716 & tmp9717) | (tmp9716 & tmp9718) | (tmp9717 & tmp9718);
  wire tmp9720;
  assign tmp9720 = 1'b0;
  wire tmp9721;
  assign tmp9721 = 1'b0;
  wire tmp9722;
  assign tmp9722 = 1'b0;
  wire tmp9723;
  assign tmp9723 = (tmp9720 & tmp9721) | (tmp9720 & tmp9722) | (tmp9721 & tmp9722);
  wire tmp9724;
  assign tmp9724 = 1'b0;
  wire tmp9725;
  assign tmp9725 = 1'b0;
  wire tmp9726;
  assign tmp9726 = 1'b0;
  wire tmp9727;
  assign tmp9727 = (tmp9724 & tmp9725) | (tmp9724 & tmp9726) | (tmp9725 & tmp9726);
  wire tmp9728;
  assign tmp9728 = (tmp9719 & tmp9723) | (tmp9719 & tmp9727) | (tmp9723 & tmp9727);
  wire tmp9729;
  assign tmp9729 = 1'b0;
  wire tmp9730;
  assign tmp9730 = 1'b0;
  wire tmp9731;
  assign tmp9731 = 1'b0;
  wire tmp9732;
  assign tmp9732 = (tmp9729 & tmp9730) | (tmp9729 & tmp9731) | (tmp9730 & tmp9731);
  wire tmp9733;
  assign tmp9733 = 1'b0;
  wire tmp9734;
  assign tmp9734 = 1'b0;
  wire tmp9735;
  assign tmp9735 = 1'b0;
  wire tmp9736;
  assign tmp9736 = (tmp9733 & tmp9734) | (tmp9733 & tmp9735) | (tmp9734 & tmp9735);
  wire tmp9737;
  assign tmp9737 = 1'b0;
  wire tmp9738;
  assign tmp9738 = 1'b0;
  wire tmp9739;
  assign tmp9739 = 1'b0;
  wire tmp9740;
  assign tmp9740 = (tmp9737 & tmp9738) | (tmp9737 & tmp9739) | (tmp9738 & tmp9739);
  wire tmp9741;
  assign tmp9741 = (tmp9732 & tmp9736) | (tmp9732 & tmp9740) | (tmp9736 & tmp9740);
  wire tmp9742;
  assign tmp9742 = 1'b0;
  wire tmp9743;
  assign tmp9743 = 1'b0;
  wire tmp9744;
  assign tmp9744 = 1'b0;
  wire tmp9745;
  assign tmp9745 = (tmp9742 & tmp9743) | (tmp9742 & tmp9744) | (tmp9743 & tmp9744);
  wire tmp9746;
  assign tmp9746 = 1'b0;
  wire tmp9747;
  assign tmp9747 = 1'b0;
  wire tmp9748;
  assign tmp9748 = 1'b0;
  wire tmp9749;
  assign tmp9749 = (tmp9746 & tmp9747) | (tmp9746 & tmp9748) | (tmp9747 & tmp9748);
  wire tmp9750;
  assign tmp9750 = 1'b0;
  wire tmp9751;
  assign tmp9751 = 1'b0;
  wire tmp9752;
  assign tmp9752 = 1'b0;
  wire tmp9753;
  assign tmp9753 = (tmp9750 & tmp9751) | (tmp9750 & tmp9752) | (tmp9751 & tmp9752);
  wire tmp9754;
  assign tmp9754 = (tmp9745 & tmp9749) | (tmp9745 & tmp9753) | (tmp9749 & tmp9753);
  wire tmp9755;
  assign tmp9755 = (tmp9728 & tmp9741) | (tmp9728 & tmp9754) | (tmp9741 & tmp9754);
  wire tmp9756;
  assign tmp9756 = 1'b0;
  wire tmp9757;
  assign tmp9757 = 1'b0;
  wire tmp9758;
  assign tmp9758 = 1'b0;
  wire tmp9759;
  assign tmp9759 = (tmp9756 & tmp9757) | (tmp9756 & tmp9758) | (tmp9757 & tmp9758);
  wire tmp9760;
  assign tmp9760 = 1'b0;
  wire tmp9761;
  assign tmp9761 = 1'b0;
  wire tmp9762;
  assign tmp9762 = 1'b0;
  wire tmp9763;
  assign tmp9763 = (tmp9760 & tmp9761) | (tmp9760 & tmp9762) | (tmp9761 & tmp9762);
  wire tmp9764;
  assign tmp9764 = 1'b0;
  wire tmp9765;
  assign tmp9765 = 1'b0;
  wire tmp9766;
  assign tmp9766 = 1'b0;
  wire tmp9767;
  assign tmp9767 = (tmp9764 & tmp9765) | (tmp9764 & tmp9766) | (tmp9765 & tmp9766);
  wire tmp9768;
  assign tmp9768 = (tmp9759 & tmp9763) | (tmp9759 & tmp9767) | (tmp9763 & tmp9767);
  wire tmp9769;
  assign tmp9769 = 1'b0;
  wire tmp9770;
  assign tmp9770 = 1'b0;
  wire tmp9771;
  assign tmp9771 = 1'b0;
  wire tmp9772;
  assign tmp9772 = (tmp9769 & tmp9770) | (tmp9769 & tmp9771) | (tmp9770 & tmp9771);
  wire tmp9773;
  assign tmp9773 = 1'b0;
  wire tmp9774;
  assign tmp9774 = 1'b0;
  wire tmp9775;
  assign tmp9775 = 1'b0;
  wire tmp9776;
  assign tmp9776 = (tmp9773 & tmp9774) | (tmp9773 & tmp9775) | (tmp9774 & tmp9775);
  wire tmp9777;
  assign tmp9777 = 1'b0;
  wire tmp9778;
  assign tmp9778 = 1'b0;
  wire tmp9779;
  assign tmp9779 = 1'b0;
  wire tmp9780;
  assign tmp9780 = (tmp9777 & tmp9778) | (tmp9777 & tmp9779) | (tmp9778 & tmp9779);
  wire tmp9781;
  assign tmp9781 = (tmp9772 & tmp9776) | (tmp9772 & tmp9780) | (tmp9776 & tmp9780);
  wire tmp9782;
  assign tmp9782 = 1'b0;
  wire tmp9783;
  assign tmp9783 = 1'b0;
  wire tmp9784;
  assign tmp9784 = 1'b0;
  wire tmp9785;
  assign tmp9785 = (tmp9782 & tmp9783) | (tmp9782 & tmp9784) | (tmp9783 & tmp9784);
  wire tmp9786;
  assign tmp9786 = 1'b0;
  wire tmp9787;
  assign tmp9787 = 1'b0;
  wire tmp9788;
  assign tmp9788 = 1'b0;
  wire tmp9789;
  assign tmp9789 = (tmp9786 & tmp9787) | (tmp9786 & tmp9788) | (tmp9787 & tmp9788);
  wire tmp9790;
  assign tmp9790 = 1'b0;
  wire tmp9791;
  assign tmp9791 = 1'b0;
  wire tmp9792;
  assign tmp9792 = 1'b0;
  wire tmp9793;
  assign tmp9793 = (tmp9790 & tmp9791) | (tmp9790 & tmp9792) | (tmp9791 & tmp9792);
  wire tmp9794;
  assign tmp9794 = (tmp9785 & tmp9789) | (tmp9785 & tmp9793) | (tmp9789 & tmp9793);
  wire tmp9795;
  assign tmp9795 = (tmp9768 & tmp9781) | (tmp9768 & tmp9794) | (tmp9781 & tmp9794);
  wire tmp9796;
  assign tmp9796 = 1'b0;
  wire tmp9797;
  assign tmp9797 = 1'b0;
  wire tmp9798;
  assign tmp9798 = 1'b0;
  wire tmp9799;
  assign tmp9799 = (tmp9796 & tmp9797) | (tmp9796 & tmp9798) | (tmp9797 & tmp9798);
  wire tmp9800;
  assign tmp9800 = 1'b0;
  wire tmp9801;
  assign tmp9801 = 1'b0;
  wire tmp9802;
  assign tmp9802 = 1'b0;
  wire tmp9803;
  assign tmp9803 = (tmp9800 & tmp9801) | (tmp9800 & tmp9802) | (tmp9801 & tmp9802);
  wire tmp9804;
  assign tmp9804 = 1'b0;
  wire tmp9805;
  assign tmp9805 = 1'b0;
  wire tmp9806;
  assign tmp9806 = 1'b0;
  wire tmp9807;
  assign tmp9807 = (tmp9804 & tmp9805) | (tmp9804 & tmp9806) | (tmp9805 & tmp9806);
  wire tmp9808;
  assign tmp9808 = (tmp9799 & tmp9803) | (tmp9799 & tmp9807) | (tmp9803 & tmp9807);
  wire tmp9809;
  assign tmp9809 = 1'b0;
  wire tmp9810;
  assign tmp9810 = 1'b0;
  wire tmp9811;
  assign tmp9811 = 1'b0;
  wire tmp9812;
  assign tmp9812 = (tmp9809 & tmp9810) | (tmp9809 & tmp9811) | (tmp9810 & tmp9811);
  wire tmp9813;
  assign tmp9813 = 1'b0;
  wire tmp9814;
  assign tmp9814 = 1'b0;
  wire tmp9815;
  assign tmp9815 = 1'b0;
  wire tmp9816;
  assign tmp9816 = (tmp9813 & tmp9814) | (tmp9813 & tmp9815) | (tmp9814 & tmp9815);
  wire tmp9817;
  assign tmp9817 = 1'b0;
  wire tmp9818;
  assign tmp9818 = 1'b0;
  wire tmp9819;
  assign tmp9819 = 1'b0;
  wire tmp9820;
  assign tmp9820 = (tmp9817 & tmp9818) | (tmp9817 & tmp9819) | (tmp9818 & tmp9819);
  wire tmp9821;
  assign tmp9821 = (tmp9812 & tmp9816) | (tmp9812 & tmp9820) | (tmp9816 & tmp9820);
  wire tmp9822;
  assign tmp9822 = 1'b0;
  wire tmp9823;
  assign tmp9823 = 1'b0;
  wire tmp9824;
  assign tmp9824 = 1'b0;
  wire tmp9825;
  assign tmp9825 = (tmp9822 & tmp9823) | (tmp9822 & tmp9824) | (tmp9823 & tmp9824);
  wire tmp9826;
  assign tmp9826 = 1'b0;
  wire tmp9827;
  assign tmp9827 = 1'b0;
  wire tmp9828;
  assign tmp9828 = 1'b0;
  wire tmp9829;
  assign tmp9829 = (tmp9826 & tmp9827) | (tmp9826 & tmp9828) | (tmp9827 & tmp9828);
  wire tmp9830;
  assign tmp9830 = 1'b0;
  wire tmp9831;
  assign tmp9831 = 1'b0;
  wire tmp9832;
  assign tmp9832 = 1'b0;
  wire tmp9833;
  assign tmp9833 = (tmp9830 & tmp9831) | (tmp9830 & tmp9832) | (tmp9831 & tmp9832);
  wire tmp9834;
  assign tmp9834 = (tmp9825 & tmp9829) | (tmp9825 & tmp9833) | (tmp9829 & tmp9833);
  wire tmp9835;
  assign tmp9835 = (tmp9808 & tmp9821) | (tmp9808 & tmp9834) | (tmp9821 & tmp9834);
  wire tmp9836;
  assign tmp9836 = (tmp9755 & tmp9795) | (tmp9755 & tmp9835) | (tmp9795 & tmp9835);
  wire tmp9837;
  assign tmp9837 = (tmp9594 & tmp9715) | (tmp9594 & tmp9836) | (tmp9715 & tmp9836);
  wire tmp9838;
  assign tmp9838 = (tmp9109 & tmp9473) | (tmp9109 & tmp9837) | (tmp9473 & tmp9837);
  wire tmp9839;
  assign tmp9839 = (tmp7652 & tmp8745) | (tmp7652 & tmp9838) | (tmp8745 & tmp9838);
  wire tmp9840;
  assign tmp9840 = (tmp3279 & tmp6559) | (tmp3279 & tmp9839) | (tmp6559 & tmp9839);
  assign po0 = tmp9840;
endmodule // test_inv
